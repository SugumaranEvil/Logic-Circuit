<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-85.0917,-33.9386,201.41,-181.701</PageViewport>
<gate>
<ID>2</ID>
<type>AA_LABEL</type>
<position>48.5,-55.5</position>
<gparam>LABEL_TEXT Half Adder</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>3</ID>
<type>AA_LABEL</type>
<position>47.5,-102.5</position>
<gparam>LABEL_TEXT Full Adder</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>4</ID>
<type>AA_LABEL</type>
<position>86.5,-128.5</position>
<gparam>LABEL_TEXT Carry</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>32</ID>
<type>GA_LED</type>
<position>74,-67.5</position>
<input>
<ID>N_in0</ID>72 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>38</ID>
<type>AA_LABEL</type>
<position>75,-63.5</position>
<gparam>LABEL_TEXT Output 0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>99</ID>
<type>AI_XOR2</type>
<position>46.5,-67.5</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>72 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>101</ID>
<type>AA_AND2</type>
<position>50.5,-76.5</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>3 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>115</ID>
<type>AA_TOGGLE</type>
<position>21,-66</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>116</ID>
<type>AA_LABEL</type>
<position>21.5,-62</position>
<gparam>LABEL_TEXT A1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>118</ID>
<type>AA_TOGGLE</type>
<position>21,-69</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>119</ID>
<type>AA_LABEL</type>
<position>21,-72</position>
<gparam>LABEL_TEXT B1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>122</ID>
<type>GA_LED</type>
<position>74,-76.5</position>
<input>
<ID>N_in0</ID>3 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>123</ID>
<type>AA_LABEL</type>
<position>75,-72.5</position>
<gparam>LABEL_TEXT Carry</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>151</ID>
<type>AI_XOR2</type>
<position>47.5,-115.5</position>
<input>
<ID>IN_0</ID>99 </input>
<input>
<ID>IN_1</ID>93 </input>
<output>
<ID>OUT</ID>94 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>153</ID>
<type>AI_XOR2</type>
<position>57.5,-125</position>
<input>
<ID>IN_0</ID>94 </input>
<input>
<ID>IN_1</ID>95 </input>
<output>
<ID>OUT</ID>96 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>155</ID>
<type>AA_TOGGLE</type>
<position>17,-114.5</position>
<output>
<ID>OUT_0</ID>99 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>157</ID>
<type>AA_TOGGLE</type>
<position>16.5,-120.5</position>
<output>
<ID>OUT_0</ID>93 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>159</ID>
<type>AA_TOGGLE</type>
<position>18,-132.5</position>
<output>
<ID>OUT_0</ID>95 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>161</ID>
<type>GA_LED</type>
<position>84,-122.5</position>
<input>
<ID>N_in0</ID>96 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>165</ID>
<type>AA_LABEL</type>
<position>18,-110.5</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>166</ID>
<type>AA_LABEL</type>
<position>17,-117.5</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>167</ID>
<type>AA_LABEL</type>
<position>18.5,-128</position>
<gparam>LABEL_TEXT C</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>168</ID>
<type>AA_LABEL</type>
<position>85,-118.5</position>
<gparam>LABEL_TEXT Output</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>170</ID>
<type>GA_LED</type>
<position>85.5,-132.5</position>
<input>
<ID>N_in0</ID>107 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>174</ID>
<type>AA_AND2</type>
<position>50,-131.5</position>
<input>
<ID>IN_0</ID>93 </input>
<input>
<ID>IN_1</ID>95 </input>
<output>
<ID>OUT</ID>106 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>176</ID>
<type>AE_OR2</type>
<position>50.5,-139</position>
<input>
<ID>IN_0</ID>93 </input>
<input>
<ID>IN_1</ID>95 </input>
<output>
<ID>OUT</ID>104 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>178</ID>
<type>AA_AND2</type>
<position>64.5,-138</position>
<input>
<ID>IN_0</ID>99 </input>
<input>
<ID>IN_1</ID>104 </input>
<output>
<ID>OUT</ID>105 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>180</ID>
<type>AE_OR2</type>
<position>75.5,-133.5</position>
<input>
<ID>IN_0</ID>106 </input>
<input>
<ID>IN_1</ID>105 </input>
<output>
<ID>OUT</ID>107 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33,-66.5,33,-66</points>
<intersection>-66.5 1</intersection>
<intersection>-66 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>33,-66.5,43.5,-66.5</points>
<connection>
<GID>99</GID>
<name>IN_0</name></connection>
<intersection>33 0</intersection>
<intersection>41.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>23,-66,33,-66</points>
<connection>
<GID>115</GID>
<name>OUT_0</name></connection>
<intersection>33 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>41.5,-75.5,41.5,-66.5</points>
<intersection>-75.5 4</intersection>
<intersection>-66.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>41.5,-75.5,47.5,-75.5</points>
<connection>
<GID>101</GID>
<name>IN_0</name></connection>
<intersection>41.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33,-69,33,-68.5</points>
<intersection>-69 2</intersection>
<intersection>-68.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>33,-68.5,43.5,-68.5</points>
<connection>
<GID>99</GID>
<name>IN_1</name></connection>
<intersection>33 0</intersection>
<intersection>37 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>23,-69,33,-69</points>
<connection>
<GID>118</GID>
<name>OUT_0</name></connection>
<intersection>33 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>37,-77.5,37,-68.5</points>
<intersection>-77.5 4</intersection>
<intersection>-68.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>37,-77.5,47.5,-77.5</points>
<connection>
<GID>101</GID>
<name>IN_1</name></connection>
<intersection>37 3</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53.5,-76.5,73,-76.5</points>
<connection>
<GID>101</GID>
<name>OUT</name></connection>
<connection>
<GID>122</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>72</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>49.5,-67.5,73,-67.5</points>
<connection>
<GID>32</GID>
<name>N_in0</name></connection>
<connection>
<GID>99</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>93</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31.5,-120.5,31.5,-116.5</points>
<intersection>-120.5 2</intersection>
<intersection>-116.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>31.5,-116.5,44.5,-116.5</points>
<connection>
<GID>151</GID>
<name>IN_1</name></connection>
<intersection>31.5 0</intersection>
<intersection>43.5 7</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>18.5,-120.5,31.5,-120.5</points>
<connection>
<GID>157</GID>
<name>OUT_0</name></connection>
<intersection>31.5 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>43.5,-130.5,43.5,-116.5</points>
<intersection>-130.5 8</intersection>
<intersection>-116.5 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>43.5,-130.5,47,-130.5</points>
<connection>
<GID>174</GID>
<name>IN_0</name></connection>
<intersection>43.5 7</intersection>
<intersection>46 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>46,-138,46,-130.5</points>
<intersection>-138 10</intersection>
<intersection>-130.5 8</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>46,-138,47.5,-138</points>
<connection>
<GID>176</GID>
<name>IN_0</name></connection>
<intersection>46 9</intersection></hsegment></shape></wire>
<wire>
<ID>94</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52.5,-124,52.5,-115.5</points>
<intersection>-124 1</intersection>
<intersection>-115.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>52.5,-124,54.5,-124</points>
<connection>
<GID>153</GID>
<name>IN_0</name></connection>
<intersection>52.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>50.5,-115.5,52.5,-115.5</points>
<connection>
<GID>151</GID>
<name>OUT</name></connection>
<intersection>52.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>95</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37,-132.5,37,-126</points>
<intersection>-132.5 2</intersection>
<intersection>-126 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>37,-126,54.5,-126</points>
<connection>
<GID>153</GID>
<name>IN_1</name></connection>
<intersection>37 0</intersection>
<intersection>42 7</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>20,-132.5,37,-132.5</points>
<connection>
<GID>159</GID>
<name>OUT_0</name></connection>
<intersection>37 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>42,-132.5,42,-126</points>
<intersection>-132.5 8</intersection>
<intersection>-126 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>42,-132.5,47,-132.5</points>
<connection>
<GID>174</GID>
<name>IN_1</name></connection>
<intersection>42 7</intersection>
<intersection>44 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>44,-140,44,-132.5</points>
<intersection>-140 10</intersection>
<intersection>-132.5 8</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>44,-140,47.5,-140</points>
<connection>
<GID>176</GID>
<name>IN_1</name></connection>
<intersection>44 9</intersection></hsegment></shape></wire>
<wire>
<ID>96</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>71.5,-125,71.5,-122.5</points>
<intersection>-125 2</intersection>
<intersection>-122.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>71.5,-122.5,83,-122.5</points>
<connection>
<GID>161</GID>
<name>N_in0</name></connection>
<intersection>71.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>60.5,-125,71.5,-125</points>
<connection>
<GID>153</GID>
<name>OUT</name></connection>
<intersection>71.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>99</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19,-114.5,44.5,-114.5</points>
<connection>
<GID>151</GID>
<name>IN_0</name></connection>
<connection>
<GID>155</GID>
<name>OUT_0</name></connection>
<intersection>41 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>41,-137,41,-114.5</points>
<intersection>-137 3</intersection>
<intersection>-114.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>41,-137,61.5,-137</points>
<connection>
<GID>178</GID>
<name>IN_0</name></connection>
<intersection>41 2</intersection></hsegment></shape></wire>
<wire>
<ID>104</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53.5,-139,61.5,-139</points>
<connection>
<GID>176</GID>
<name>OUT</name></connection>
<connection>
<GID>178</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>105</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>69.5,-138,69.5,-134.5</points>
<intersection>-138 2</intersection>
<intersection>-134.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>69.5,-134.5,72.5,-134.5</points>
<connection>
<GID>180</GID>
<name>IN_1</name></connection>
<intersection>69.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>67.5,-138,69.5,-138</points>
<connection>
<GID>178</GID>
<name>OUT</name></connection>
<intersection>69.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>106</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>62.5,-132.5,62.5,-131.5</points>
<intersection>-132.5 1</intersection>
<intersection>-131.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>62.5,-132.5,72.5,-132.5</points>
<connection>
<GID>180</GID>
<name>IN_0</name></connection>
<intersection>62.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>53,-131.5,62.5,-131.5</points>
<connection>
<GID>174</GID>
<name>OUT</name></connection>
<intersection>62.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>107</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>81.5,-133.5,81.5,-132.5</points>
<intersection>-133.5 2</intersection>
<intersection>-132.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>81.5,-132.5,84.5,-132.5</points>
<connection>
<GID>170</GID>
<name>N_in0</name></connection>
<intersection>81.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>78.5,-133.5,81.5,-133.5</points>
<connection>
<GID>180</GID>
<name>OUT</name></connection>
<intersection>81.5 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,3.46927e-006,177.8,-91.7</PageViewport></page 1>
<page 2>
<PageViewport>0,3.46927e-006,177.8,-91.7</PageViewport></page 2>
<page 3>
<PageViewport>0,3.46927e-006,177.8,-91.7</PageViewport></page 3>
<page 4>
<PageViewport>0,3.46927e-006,177.8,-91.7</PageViewport></page 4>
<page 5>
<PageViewport>0,3.46927e-006,177.8,-91.7</PageViewport></page 5>
<page 6>
<PageViewport>0,3.46927e-006,177.8,-91.7</PageViewport></page 6>
<page 7>
<PageViewport>0,3.46927e-006,177.8,-91.7</PageViewport></page 7>
<page 8>
<PageViewport>0,3.46927e-006,177.8,-91.7</PageViewport></page 8>
<page 9>
<PageViewport>0,3.46927e-006,177.8,-91.7</PageViewport></page 9></circuit>