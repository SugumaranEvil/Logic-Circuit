<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-78.23,-21.4136,176.438,-152.758</PageViewport>
<gate>
<ID>1</ID>
<type>AA_LABEL</type>
<position>45,-35.5</position>
<gparam>LABEL_TEXT Half Subtractor</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2</ID>
<type>GA_LED</type>
<position>59.5,-47.5</position>
<input>
<ID>N_in0</ID>4 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>3</ID>
<type>AA_LABEL</type>
<position>62,-44</position>
<gparam>LABEL_TEXT Output </gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>4</ID>
<type>AI_XOR2</type>
<position>43,-47.5</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>4 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5</ID>
<type>AA_AND2</type>
<position>53,-56.5</position>
<input>
<ID>IN_0</ID>6 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>3 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_TOGGLE</type>
<position>17.5,-46</position>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>7</ID>
<type>AA_LABEL</type>
<position>18,-42</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>8</ID>
<type>AA_TOGGLE</type>
<position>17.5,-49</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>9</ID>
<type>AA_LABEL</type>
<position>17.5,-52</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>10</ID>
<type>GA_LED</type>
<position>66.5,-56.5</position>
<input>
<ID>N_in0</ID>3 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>11</ID>
<type>AA_LABEL</type>
<position>67.5,-53</position>
<gparam>LABEL_TEXT Borrow</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>12</ID>
<type>AI_XOR2</type>
<position>27,-87.5</position>
<input>
<ID>IN_0</ID>12 </input>
<input>
<ID>IN_1</ID>13 </input>
<output>
<ID>OUT</ID>15 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>13</ID>
<type>AA_INVERTER</type>
<position>43.5,-54.5</position>
<input>
<ID>IN_0</ID>5 </input>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>14</ID>
<type>AA_AND2</type>
<position>35,-102.5</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>13 </input>
<output>
<ID>OUT</ID>10 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>15</ID>
<type>AA_INVERTER</type>
<position>28.5,-101.5</position>
<input>
<ID>IN_0</ID>12 </input>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>16</ID>
<type>AI_XOR2</type>
<position>47.5,-88.5</position>
<input>
<ID>IN_0</ID>15 </input>
<input>
<ID>IN_1</ID>11 </input>
<output>
<ID>OUT</ID>16 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>17</ID>
<type>AA_AND2</type>
<position>54,-97</position>
<input>
<ID>IN_0</ID>7 </input>
<input>
<ID>IN_1</ID>11 </input>
<output>
<ID>OUT</ID>9 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>18</ID>
<type>AA_INVERTER</type>
<position>47.5,-96</position>
<input>
<ID>IN_0</ID>15 </input>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>19</ID>
<type>AE_OR2</type>
<position>65,-99</position>
<input>
<ID>IN_0</ID>9 </input>
<input>
<ID>IN_1</ID>10 </input>
<output>
<ID>OUT</ID>14 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>20</ID>
<type>GA_LED</type>
<position>75,-99</position>
<input>
<ID>N_in0</ID>14 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>21</ID>
<type>AA_TOGGLE</type>
<position>-2.5,-86.5</position>
<output>
<ID>OUT_0</ID>12 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>22</ID>
<type>AA_LABEL</type>
<position>-2.5,-82.5</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>23</ID>
<type>AA_TOGGLE</type>
<position>-2.5,-90</position>
<output>
<ID>OUT_0</ID>13 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>24</ID>
<type>AA_LABEL</type>
<position>-2.5,-92.5</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>25</ID>
<type>AA_TOGGLE</type>
<position>-2,-98</position>
<output>
<ID>OUT_0</ID>11 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>26</ID>
<type>AA_LABEL</type>
<position>-2.5,-100.5</position>
<gparam>LABEL_TEXT C</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>27</ID>
<type>GA_LED</type>
<position>71.5,-88.5</position>
<input>
<ID>N_in0</ID>16 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>28</ID>
<type>AA_LABEL</type>
<position>37.5,-76.5</position>
<gparam>LABEL_TEXT Full Subtractor</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>29</ID>
<type>AA_LABEL</type>
<position>70.5,-84</position>
<gparam>LABEL_TEXT Output </gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>30</ID>
<type>AA_LABEL</type>
<position>74,-95.5</position>
<gparam>LABEL_TEXT Borrow</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>31.5,-101.5,32,-101.5</points>
<connection>
<GID>14</GID>
<name>IN_0</name></connection>
<connection>
<GID>15</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29.5,-49,29.5,-48.5</points>
<intersection>-49 2</intersection>
<intersection>-48.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29.5,-48.5,40,-48.5</points>
<connection>
<GID>4</GID>
<name>IN_1</name></connection>
<intersection>29.5 0</intersection>
<intersection>33.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>19.5,-49,29.5,-49</points>
<connection>
<GID>8</GID>
<name>OUT_0</name></connection>
<intersection>29.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>33.5,-57.5,33.5,-48.5</points>
<intersection>-57.5 4</intersection>
<intersection>-48.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>33.5,-57.5,50,-57.5</points>
<connection>
<GID>5</GID>
<name>IN_1</name></connection>
<intersection>33.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>56,-56.5,65.5,-56.5</points>
<connection>
<GID>5</GID>
<name>OUT</name></connection>
<connection>
<GID>10</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<hsegment>
<ID>10</ID>
<points>46,-47.5,58.5,-47.5</points>
<connection>
<GID>2</GID>
<name>N_in0</name></connection>
<connection>
<GID>4</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37.5,-54.5,37.5,-46</points>
<intersection>-54.5 1</intersection>
<intersection>-46.5 2</intersection>
<intersection>-46 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>37.5,-54.5,40.5,-54.5</points>
<connection>
<GID>13</GID>
<name>IN_0</name></connection>
<intersection>37.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>37.5,-46.5,40,-46.5</points>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<intersection>37.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>19.5,-46,37.5,-46</points>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<intersection>37.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>48,-55.5,48,-54.5</points>
<intersection>-55.5 1</intersection>
<intersection>-54.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>48,-55.5,50,-55.5</points>
<connection>
<GID>5</GID>
<name>IN_0</name></connection>
<intersection>48 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>46.5,-54.5,48,-54.5</points>
<connection>
<GID>13</GID>
<name>OUT_0</name></connection>
<intersection>48 0</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>50.5,-96,51,-96</points>
<connection>
<GID>17</GID>
<name>IN_0</name></connection>
<connection>
<GID>18</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>59.5,-98,59.5,-97</points>
<intersection>-98 1</intersection>
<intersection>-97 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>59.5,-98,62,-98</points>
<connection>
<GID>19</GID>
<name>IN_0</name></connection>
<intersection>59.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>57,-97,59.5,-97</points>
<connection>
<GID>17</GID>
<name>OUT</name></connection>
<intersection>59.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50,-102.5,50,-100</points>
<intersection>-102.5 2</intersection>
<intersection>-100 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50,-100,62,-100</points>
<connection>
<GID>19</GID>
<name>IN_1</name></connection>
<intersection>50 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>38,-102.5,50,-102.5</points>
<connection>
<GID>14</GID>
<name>OUT</name></connection>
<intersection>50 0</intersection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>2</ID>
<points>41.5,-98,41.5,-89.5</points>
<intersection>-98 3</intersection>
<intersection>-89.5 4</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>0,-98,51,-98</points>
<connection>
<GID>17</GID>
<name>IN_1</name></connection>
<connection>
<GID>25</GID>
<name>OUT_0</name></connection>
<intersection>41.5 2</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>41.5,-89.5,44.5,-89.5</points>
<connection>
<GID>16</GID>
<name>IN_1</name></connection>
<intersection>41.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-0.5,-86.5,24,-86.5</points>
<connection>
<GID>12</GID>
<name>IN_0</name></connection>
<connection>
<GID>21</GID>
<name>OUT_0</name></connection>
<intersection>22.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>22.5,-101.5,22.5,-86.5</points>
<intersection>-101.5 4</intersection>
<intersection>-86.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>22.5,-101.5,25.5,-101.5</points>
<connection>
<GID>15</GID>
<name>IN_0</name></connection>
<intersection>22.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>20.5,-88.5,24,-88.5</points>
<connection>
<GID>12</GID>
<name>IN_1</name></connection>
<intersection>20.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>20.5,-103.5,20.5,-88.5</points>
<intersection>-103.5 4</intersection>
<intersection>-90 5</intersection>
<intersection>-88.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>20.5,-103.5,32,-103.5</points>
<connection>
<GID>14</GID>
<name>IN_1</name></connection>
<intersection>20.5 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-0.5,-90,20.5,-90</points>
<connection>
<GID>23</GID>
<name>OUT_0</name></connection>
<intersection>20.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>68,-99,74,-99</points>
<connection>
<GID>19</GID>
<name>OUT</name></connection>
<connection>
<GID>20</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>30,-87.5,44.5,-87.5</points>
<connection>
<GID>16</GID>
<name>IN_0</name></connection>
<connection>
<GID>12</GID>
<name>OUT</name></connection>
<intersection>38 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>38,-96,38,-87.5</points>
<intersection>-96 4</intersection>
<intersection>-87.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>38,-96,44.5,-96</points>
<connection>
<GID>18</GID>
<name>IN_0</name></connection>
<intersection>38 3</intersection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>50.5,-88.5,70.5,-88.5</points>
<connection>
<GID>16</GID>
<name>OUT</name></connection>
<connection>
<GID>27</GID>
<name>N_in0</name></connection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,4.48114e-006,177.8,-91.7</PageViewport></page 1>
<page 2>
<PageViewport>0,4.48114e-006,177.8,-91.7</PageViewport></page 2>
<page 3>
<PageViewport>0,4.48114e-006,177.8,-91.7</PageViewport></page 3>
<page 4>
<PageViewport>0,4.48114e-006,177.8,-91.7</PageViewport></page 4>
<page 5>
<PageViewport>0,4.48114e-006,177.8,-91.7</PageViewport></page 5>
<page 6>
<PageViewport>0,4.48114e-006,177.8,-91.7</PageViewport></page 6>
<page 7>
<PageViewport>0,4.48114e-006,177.8,-91.7</PageViewport></page 7>
<page 8>
<PageViewport>0,4.48114e-006,177.8,-91.7</PageViewport></page 8>
<page 9>
<PageViewport>0,4.48114e-006,177.8,-91.7</PageViewport></page 9></circuit>