<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-145.686,-104.039,363.652,-366.729</PageViewport>
<gate>
<ID>1</ID>
<type>AI_XOR2</type>
<position>32.5,-138.5</position>
<input>
<ID>IN_0</ID>31 </input>
<input>
<ID>IN_1</ID>30 </input>
<output>
<ID>OUT</ID>18 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>11</ID>
<type>GA_LED</type>
<position>89,-138.5</position>
<input>
<ID>N_in0</ID>18 </input>
<input>
<ID>N_in1</ID>100 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>13</ID>
<type>AA_LABEL</type>
<position>-12,-134.5</position>
<gparam>LABEL_TEXT A0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>16</ID>
<type>AA_LABEL</type>
<position>-2.5,-141</position>
<gparam>LABEL_TEXT B0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>18</ID>
<type>AA_LABEL</type>
<position>-10.5,-150</position>
<gparam>LABEL_TEXT A1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>32</ID>
<type>AA_LABEL</type>
<position>90,-135</position>
<gparam>LABEL_TEXT Output BIT 0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>35</ID>
<type>GA_LED</type>
<position>67.5,-166</position>
<input>
<ID>N_in0</ID>17 </input>
<input>
<ID>N_in1</ID>96 </input>
<input>
<ID>N_in2</ID>96 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>36</ID>
<type>AA_AND2</type>
<position>40.5,-165</position>
<input>
<ID>IN_0</ID>32 </input>
<input>
<ID>IN_1</ID>21 </input>
<output>
<ID>OUT</ID>16 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>37</ID>
<type>AE_OR2</type>
<position>40.5,-171.5</position>
<input>
<ID>IN_0</ID>32 </input>
<input>
<ID>IN_1</ID>21 </input>
<output>
<ID>OUT</ID>14 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>38</ID>
<type>AA_AND2</type>
<position>49.5,-170.5</position>
<input>
<ID>IN_0</ID>19 </input>
<input>
<ID>IN_1</ID>14 </input>
<output>
<ID>OUT</ID>15 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>39</ID>
<type>AE_OR2</type>
<position>60.5,-166</position>
<input>
<ID>IN_0</ID>16 </input>
<input>
<ID>IN_1</ID>15 </input>
<output>
<ID>OUT</ID>17 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>41</ID>
<type>AA_AND2</type>
<position>38.5,-146.5</position>
<input>
<ID>IN_0</ID>31 </input>
<input>
<ID>IN_1</ID>30 </input>
<output>
<ID>OUT</ID>19 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>43</ID>
<type>AA_LABEL</type>
<position>-2.5,-156</position>
<gparam>LABEL_TEXT B1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>45</ID>
<type>AI_XOR2</type>
<position>46.5,-151</position>
<input>
<ID>IN_0</ID>19 </input>
<input>
<ID>IN_1</ID>32 </input>
<output>
<ID>OUT</ID>20 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>47</ID>
<type>AI_XOR2</type>
<position>59,-156.5</position>
<input>
<ID>IN_0</ID>20 </input>
<input>
<ID>IN_1</ID>21 </input>
<output>
<ID>OUT</ID>22 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>48</ID>
<type>GA_LED</type>
<position>89.5,-156.5</position>
<input>
<ID>N_in0</ID>22 </input>
<input>
<ID>N_in1</ID>101 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>49</ID>
<type>AA_LABEL</type>
<position>90.5,-153</position>
<gparam>LABEL_TEXT Output BIT1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>62</ID>
<type>AA_LABEL</type>
<position>-9,-179.5</position>
<gparam>LABEL_TEXT A2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>63</ID>
<type>GA_LED</type>
<position>67.5,-195</position>
<input>
<ID>N_in0</ID>36 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>64</ID>
<type>AA_AND2</type>
<position>40,-194</position>
<input>
<ID>IN_0</ID>41 </input>
<input>
<ID>IN_1</ID>39 </input>
<output>
<ID>OUT</ID>35 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>65</ID>
<type>AE_OR2</type>
<position>40,-200.5</position>
<input>
<ID>IN_0</ID>41 </input>
<input>
<ID>IN_1</ID>39 </input>
<output>
<ID>OUT</ID>33 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>66</ID>
<type>AA_AND2</type>
<position>49,-199.5</position>
<input>
<ID>IN_0</ID>17 </input>
<input>
<ID>IN_1</ID>33 </input>
<output>
<ID>OUT</ID>34 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>67</ID>
<type>AE_OR2</type>
<position>60,-195</position>
<input>
<ID>IN_0</ID>35 </input>
<input>
<ID>IN_1</ID>34 </input>
<output>
<ID>OUT</ID>36 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>69</ID>
<type>AA_LABEL</type>
<position>-2.5,-184.5</position>
<gparam>LABEL_TEXT B2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>70</ID>
<type>AI_XOR2</type>
<position>46,-180</position>
<input>
<ID>IN_0</ID>17 </input>
<input>
<ID>IN_1</ID>41 </input>
<output>
<ID>OUT</ID>38 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>71</ID>
<type>AI_XOR2</type>
<position>58.5,-185.5</position>
<input>
<ID>IN_0</ID>38 </input>
<input>
<ID>IN_1</ID>39 </input>
<output>
<ID>OUT</ID>40 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>72</ID>
<type>GA_LED</type>
<position>90,-185.5</position>
<input>
<ID>N_in0</ID>40 </input>
<input>
<ID>N_in1</ID>102 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>73</ID>
<type>AA_LABEL</type>
<position>91,-182</position>
<gparam>LABEL_TEXT Output BIT 2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>75</ID>
<type>AA_LABEL</type>
<position>-8,-207.5</position>
<gparam>LABEL_TEXT A3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>76</ID>
<type>GA_LED</type>
<position>69.5,-222.5</position>
<input>
<ID>N_in0</ID>51 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>77</ID>
<type>AA_AND2</type>
<position>39.5,-222.5</position>
<input>
<ID>IN_0</ID>50 </input>
<input>
<ID>IN_1</ID>48 </input>
<output>
<ID>OUT</ID>45 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>78</ID>
<type>AE_OR2</type>
<position>39.5,-229</position>
<input>
<ID>IN_0</ID>50 </input>
<input>
<ID>IN_1</ID>48 </input>
<output>
<ID>OUT</ID>43 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>79</ID>
<type>AA_AND2</type>
<position>48.5,-228</position>
<input>
<ID>IN_0</ID>36 </input>
<input>
<ID>IN_1</ID>43 </input>
<output>
<ID>OUT</ID>44 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>80</ID>
<type>AE_OR2</type>
<position>59.5,-223.5</position>
<input>
<ID>IN_0</ID>45 </input>
<input>
<ID>IN_1</ID>44 </input>
<output>
<ID>OUT</ID>51 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>82</ID>
<type>AA_LABEL</type>
<position>-1.5,-213</position>
<gparam>LABEL_TEXT B3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>83</ID>
<type>AI_XOR2</type>
<position>45.5,-208.5</position>
<input>
<ID>IN_0</ID>36 </input>
<input>
<ID>IN_1</ID>50 </input>
<output>
<ID>OUT</ID>47 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>84</ID>
<type>AI_XOR2</type>
<position>58,-214</position>
<input>
<ID>IN_0</ID>47 </input>
<input>
<ID>IN_1</ID>48 </input>
<output>
<ID>OUT</ID>49 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>85</ID>
<type>GA_LED</type>
<position>90,-214</position>
<input>
<ID>N_in0</ID>49 </input>
<input>
<ID>N_in1</ID>103 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>86</ID>
<type>AA_LABEL</type>
<position>91,-210.5</position>
<gparam>LABEL_TEXT Output BIT 3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>88</ID>
<type>AA_LABEL</type>
<position>-6.5,-237.5</position>
<gparam>LABEL_TEXT A4</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>89</ID>
<type>GA_LED</type>
<position>69.5,-252.5</position>
<input>
<ID>N_in0</ID>60 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>90</ID>
<type>AA_AND2</type>
<position>39.5,-252.5</position>
<input>
<ID>IN_0</ID>59 </input>
<input>
<ID>IN_1</ID>57 </input>
<output>
<ID>OUT</ID>54 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>91</ID>
<type>AE_OR2</type>
<position>39.5,-259</position>
<input>
<ID>IN_0</ID>59 </input>
<input>
<ID>IN_1</ID>57 </input>
<output>
<ID>OUT</ID>52 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>92</ID>
<type>AA_AND2</type>
<position>48.5,-258</position>
<input>
<ID>IN_0</ID>51 </input>
<input>
<ID>IN_1</ID>52 </input>
<output>
<ID>OUT</ID>53 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>93</ID>
<type>AE_OR2</type>
<position>59.5,-253.5</position>
<input>
<ID>IN_0</ID>54 </input>
<input>
<ID>IN_1</ID>53 </input>
<output>
<ID>OUT</ID>60 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>95</ID>
<type>AA_LABEL</type>
<position>1,-243</position>
<gparam>LABEL_TEXT B4</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>96</ID>
<type>AI_XOR2</type>
<position>45.5,-238.5</position>
<input>
<ID>IN_0</ID>51 </input>
<input>
<ID>IN_1</ID>59 </input>
<output>
<ID>OUT</ID>56 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>97</ID>
<type>AI_XOR2</type>
<position>58,-244</position>
<input>
<ID>IN_0</ID>56 </input>
<input>
<ID>IN_1</ID>57 </input>
<output>
<ID>OUT</ID>58 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>98</ID>
<type>GA_LED</type>
<position>89.5,-244</position>
<input>
<ID>N_in0</ID>58 </input>
<input>
<ID>N_in1</ID>104 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>99</ID>
<type>AA_LABEL</type>
<position>90.5,-240.5</position>
<gparam>LABEL_TEXT Output BIT 4</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>101</ID>
<type>AA_LABEL</type>
<position>-6.5,-265.5</position>
<gparam>LABEL_TEXT A5</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>102</ID>
<type>GA_LED</type>
<position>67,-282.5</position>
<input>
<ID>N_in0</ID>69 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>103</ID>
<type>AA_AND2</type>
<position>36,-281.5</position>
<input>
<ID>IN_0</ID>68 </input>
<input>
<ID>IN_1</ID>66 </input>
<output>
<ID>OUT</ID>63 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>104</ID>
<type>AE_OR2</type>
<position>36,-288</position>
<input>
<ID>IN_0</ID>68 </input>
<input>
<ID>IN_1</ID>66 </input>
<output>
<ID>OUT</ID>61 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>105</ID>
<type>AA_AND2</type>
<position>45,-287</position>
<input>
<ID>IN_0</ID>60 </input>
<input>
<ID>IN_1</ID>61 </input>
<output>
<ID>OUT</ID>62 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>106</ID>
<type>AE_OR2</type>
<position>56,-282.5</position>
<input>
<ID>IN_0</ID>63 </input>
<input>
<ID>IN_1</ID>62 </input>
<output>
<ID>OUT</ID>69 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>108</ID>
<type>AA_LABEL</type>
<position>1.5,-272</position>
<gparam>LABEL_TEXT B5</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>109</ID>
<type>AI_XOR2</type>
<position>42,-267.5</position>
<input>
<ID>IN_0</ID>60 </input>
<input>
<ID>IN_1</ID>68 </input>
<output>
<ID>OUT</ID>65 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>110</ID>
<type>AI_XOR2</type>
<position>54.5,-273</position>
<input>
<ID>IN_0</ID>65 </input>
<input>
<ID>IN_1</ID>66 </input>
<output>
<ID>OUT</ID>67 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>111</ID>
<type>GA_LED</type>
<position>90,-273</position>
<input>
<ID>N_in0</ID>67 </input>
<input>
<ID>N_in1</ID>105 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>112</ID>
<type>AA_LABEL</type>
<position>91,-269.5</position>
<gparam>LABEL_TEXT Output BIT 5</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>114</ID>
<type>AA_LABEL</type>
<position>-6.5,-294</position>
<gparam>LABEL_TEXT A6</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>115</ID>
<type>GA_LED</type>
<position>64,-311</position>
<input>
<ID>N_in0</ID>78 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>116</ID>
<type>AA_AND2</type>
<position>34,-310</position>
<input>
<ID>IN_0</ID>77 </input>
<input>
<ID>IN_1</ID>75 </input>
<output>
<ID>OUT</ID>72 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>117</ID>
<type>AE_OR2</type>
<position>34,-316.5</position>
<input>
<ID>IN_0</ID>77 </input>
<input>
<ID>IN_1</ID>75 </input>
<output>
<ID>OUT</ID>70 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>118</ID>
<type>AA_AND2</type>
<position>43,-315.5</position>
<input>
<ID>IN_0</ID>69 </input>
<input>
<ID>IN_1</ID>70 </input>
<output>
<ID>OUT</ID>71 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>119</ID>
<type>AE_OR2</type>
<position>54,-311</position>
<input>
<ID>IN_0</ID>72 </input>
<input>
<ID>IN_1</ID>71 </input>
<output>
<ID>OUT</ID>78 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>121</ID>
<type>AA_LABEL</type>
<position>2,-300.5</position>
<gparam>LABEL_TEXT B6</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>122</ID>
<type>AI_XOR2</type>
<position>40,-296</position>
<input>
<ID>IN_0</ID>69 </input>
<input>
<ID>IN_1</ID>77 </input>
<output>
<ID>OUT</ID>74 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>123</ID>
<type>AI_XOR2</type>
<position>52.5,-301.5</position>
<input>
<ID>IN_0</ID>74 </input>
<input>
<ID>IN_1</ID>75 </input>
<output>
<ID>OUT</ID>76 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>124</ID>
<type>GA_LED</type>
<position>90,-301.5</position>
<input>
<ID>N_in0</ID>76 </input>
<input>
<ID>N_in1</ID>106 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>125</ID>
<type>AA_LABEL</type>
<position>91,-298</position>
<gparam>LABEL_TEXT Output BIT 6</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>127</ID>
<type>AA_LABEL</type>
<position>-6.5,-324</position>
<gparam>LABEL_TEXT A7</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>128</ID>
<type>GA_LED</type>
<position>78.5,-340</position>
<input>
<ID>N_in0</ID>87 </input>
<input>
<ID>N_in1</ID>99 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>129</ID>
<type>AA_AND2</type>
<position>33.5,-339</position>
<input>
<ID>IN_0</ID>86 </input>
<input>
<ID>IN_1</ID>84 </input>
<output>
<ID>OUT</ID>81 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>130</ID>
<type>AE_OR2</type>
<position>33.5,-345.5</position>
<input>
<ID>IN_0</ID>86 </input>
<input>
<ID>IN_1</ID>84 </input>
<output>
<ID>OUT</ID>79 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>131</ID>
<type>AA_AND2</type>
<position>42.5,-344.5</position>
<input>
<ID>IN_0</ID>78 </input>
<input>
<ID>IN_1</ID>79 </input>
<output>
<ID>OUT</ID>80 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>132</ID>
<type>AE_OR2</type>
<position>53.5,-340</position>
<input>
<ID>IN_0</ID>81 </input>
<input>
<ID>IN_1</ID>80 </input>
<output>
<ID>OUT</ID>87 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>134</ID>
<type>AA_LABEL</type>
<position>2,-329.5</position>
<gparam>LABEL_TEXT B7</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>135</ID>
<type>AI_XOR2</type>
<position>39.5,-325</position>
<input>
<ID>IN_0</ID>78 </input>
<input>
<ID>IN_1</ID>86 </input>
<output>
<ID>OUT</ID>83 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>136</ID>
<type>AI_XOR2</type>
<position>52,-330.5</position>
<input>
<ID>IN_0</ID>83 </input>
<input>
<ID>IN_1</ID>84 </input>
<output>
<ID>OUT</ID>85 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>137</ID>
<type>GA_LED</type>
<position>89.5,-330.5</position>
<input>
<ID>N_in0</ID>85 </input>
<input>
<ID>N_in1</ID>107 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>138</ID>
<type>AA_LABEL</type>
<position>90.5,-327</position>
<gparam>LABEL_TEXT Output BIT 7</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>153</ID>
<type>AA_LABEL</type>
<position>80,-343</position>
<gparam>LABEL_TEXT Carry</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>161</ID>
<type>DD_KEYPAD_HEX</type>
<position>-48,-175</position>
<output>
<ID>OUT_0</ID>31 </output>
<output>
<ID>OUT_1</ID>32 </output>
<output>
<ID>OUT_2</ID>41 </output>
<output>
<ID>OUT_3</ID>50 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 15</lparam></gate>
<gate>
<ID>163</ID>
<type>DD_KEYPAD_HEX</type>
<position>-48.5,-194</position>
<output>
<ID>OUT_0</ID>30 </output>
<output>
<ID>OUT_1</ID>21 </output>
<output>
<ID>OUT_2</ID>39 </output>
<output>
<ID>OUT_3</ID>48 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 15</lparam></gate>
<gate>
<ID>165</ID>
<type>DD_KEYPAD_HEX</type>
<position>-53,-278.5</position>
<output>
<ID>OUT_0</ID>59 </output>
<output>
<ID>OUT_1</ID>68 </output>
<output>
<ID>OUT_2</ID>77 </output>
<output>
<ID>OUT_3</ID>86 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 15</lparam></gate>
<gate>
<ID>167</ID>
<type>DD_KEYPAD_HEX</type>
<position>-53.5,-296.5</position>
<output>
<ID>OUT_0</ID>57 </output>
<output>
<ID>OUT_1</ID>66 </output>
<output>
<ID>OUT_2</ID>75 </output>
<output>
<ID>OUT_3</ID>84 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 15</lparam></gate>
<gate>
<ID>169</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>181,-226</position>
<input>
<ID>IN_0</ID>100 </input>
<input>
<ID>IN_1</ID>101 </input>
<input>
<ID>IN_2</ID>102 </input>
<input>
<ID>IN_3</ID>103 </input>
<input>
<ID>IN_4</ID>104 </input>
<input>
<ID>IN_5</ID>105 </input>
<input>
<ID>IN_6</ID>106 </input>
<input>
<ID>IN_7</ID>107 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 254</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>171</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>172.5,-339</position>
<input>
<ID>IN_0</ID>99 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>173</ID>
<type>AA_LABEL</type>
<position>-77.5,-176.5</position>
<gparam>LABEL_TEXT 1st number_1st 4bit</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>174</ID>
<type>AA_LABEL</type>
<position>-78,-193</position>
<gparam>LABEL_TEXT 2nd number_1st 4bit</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>175</ID>
<type>AA_LABEL</type>
<position>-81.5,-276</position>
<gparam>LABEL_TEXT 1st number_2nd 4bit</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>176</ID>
<type>AA_LABEL</type>
<position>-81.5,-295</position>
<gparam>LABEL_TEXT 2nd number_2nd 4bit</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>177</ID>
<type>AA_LABEL</type>
<position>180,-340</position>
<gparam>LABEL_TEXT Carry</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>178</ID>
<type>AA_LABEL</type>
<position>70,-310.5</position>
<gparam>LABEL_TEXT Carry</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>179</ID>
<type>AA_LABEL</type>
<position>73,-283</position>
<gparam>LABEL_TEXT Carry</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>180</ID>
<type>AA_LABEL</type>
<position>76,-253</position>
<gparam>LABEL_TEXT Carry</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>181</ID>
<type>AA_LABEL</type>
<position>77.5,-221.5</position>
<gparam>LABEL_TEXT Carry</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>182</ID>
<type>AA_LABEL</type>
<position>74.5,-195</position>
<gparam>LABEL_TEXT Carry</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>183</ID>
<type>AA_LABEL</type>
<position>75,-165</position>
<gparam>LABEL_TEXT Carry</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>185</ID>
<type>AA_LABEL</type>
<position>38.5,-120</position>
<gparam>LABEL_TEXT 8bit adder</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>187</ID>
<type>AA_LABEL</type>
<position>181.5,-212.5</position>
<gparam>LABEL_TEXT Output</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>14</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>43.5,-171.5,46.5,-171.5</points>
<connection>
<GID>37</GID>
<name>OUT</name></connection>
<connection>
<GID>38</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54.5,-170.5,54.5,-167</points>
<intersection>-170.5 2</intersection>
<intersection>-167 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>54.5,-167,57.5,-167</points>
<connection>
<GID>39</GID>
<name>IN_1</name></connection>
<intersection>54.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>52.5,-170.5,54.5,-170.5</points>
<connection>
<GID>38</GID>
<name>OUT</name></connection>
<intersection>54.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>43.5,-165,57.5,-165</points>
<connection>
<GID>36</GID>
<name>OUT</name></connection>
<connection>
<GID>39</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>63.5,-166,66.5,-166</points>
<connection>
<GID>39</GID>
<name>OUT</name></connection>
<connection>
<GID>35</GID>
<name>N_in0</name></connection>
<intersection>64 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>64,-179,64,-166</points>
<intersection>-179 5</intersection>
<intersection>-166 2</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>42.5,-179,64,-179</points>
<connection>
<GID>70</GID>
<name>IN_0</name></connection>
<intersection>42.5 7</intersection>
<intersection>64 3</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>42.5,-198.5,42.5,-179</points>
<intersection>-198.5 8</intersection>
<intersection>-179 5</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>42.5,-198.5,46,-198.5</points>
<connection>
<GID>66</GID>
<name>IN_0</name></connection>
<intersection>42.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>35.5,-138.5,88,-138.5</points>
<connection>
<GID>11</GID>
<name>N_in0</name></connection>
<connection>
<GID>1</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>42.5,-150,42.5,-146.5</points>
<intersection>-150 1</intersection>
<intersection>-146.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>42.5,-150,43.5,-150</points>
<connection>
<GID>45</GID>
<name>IN_0</name></connection>
<intersection>42.5 0</intersection>
<intersection>43 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>41.5,-146.5,42.5,-146.5</points>
<connection>
<GID>41</GID>
<name>OUT</name></connection>
<intersection>42.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>43,-169.5,43,-150</points>
<intersection>-169.5 4</intersection>
<intersection>-150 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>43,-169.5,46.5,-169.5</points>
<connection>
<GID>38</GID>
<name>IN_0</name></connection>
<intersection>43 3</intersection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52.5,-155.5,52.5,-151</points>
<intersection>-155.5 1</intersection>
<intersection>-151 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>52.5,-155.5,56,-155.5</points>
<connection>
<GID>47</GID>
<name>IN_0</name></connection>
<intersection>52.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>49.5,-151,52.5,-151</points>
<connection>
<GID>45</GID>
<name>OUT</name></connection>
<intersection>52.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-21.5,-157.5,56,-157.5</points>
<connection>
<GID>47</GID>
<name>IN_1</name></connection>
<intersection>-21.5 9</intersection>
<intersection>35.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>35.5,-172.5,35.5,-157.5</points>
<intersection>-172.5 6</intersection>
<intersection>-166 4</intersection>
<intersection>-157.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>35.5,-166,37.5,-166</points>
<connection>
<GID>36</GID>
<name>IN_1</name></connection>
<intersection>35.5 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>35.5,-172.5,37.5,-172.5</points>
<connection>
<GID>37</GID>
<name>IN_1</name></connection>
<intersection>35.5 3</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>-21.5,-195,-21.5,-157.5</points>
<intersection>-195 10</intersection>
<intersection>-157.5 1</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>-43.5,-195,-21.5,-195</points>
<connection>
<GID>163</GID>
<name>OUT_1</name></connection>
<intersection>-21.5 9</intersection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>62,-156.5,88.5,-156.5</points>
<connection>
<GID>47</GID>
<name>OUT</name></connection>
<connection>
<GID>48</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17,-143,17,-139.5</points>
<intersection>-143 2</intersection>
<intersection>-139.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>17,-139.5,29.5,-139.5</points>
<connection>
<GID>1</GID>
<name>IN_1</name></connection>
<intersection>17 0</intersection>
<intersection>28.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-18,-143,17,-143</points>
<intersection>-18 5</intersection>
<intersection>17 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>28.5,-147.5,28.5,-139.5</points>
<intersection>-147.5 4</intersection>
<intersection>-139.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>28.5,-147.5,35.5,-147.5</points>
<connection>
<GID>41</GID>
<name>IN_1</name></connection>
<intersection>28.5 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-18,-197,-18,-143</points>
<intersection>-197 6</intersection>
<intersection>-143 2</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-43.5,-197,-18,-197</points>
<connection>
<GID>163</GID>
<name>OUT_0</name></connection>
<intersection>-18 5</intersection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-39.5,-137.5,29.5,-137.5</points>
<connection>
<GID>1</GID>
<name>IN_0</name></connection>
<intersection>-39.5 16</intersection>
<intersection>26 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>26,-145.5,26,-137.5</points>
<intersection>-145.5 4</intersection>
<intersection>-137.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>26,-145.5,35.5,-145.5</points>
<connection>
<GID>41</GID>
<name>IN_0</name></connection>
<intersection>26 3</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>-39.5,-178,-39.5,-137.5</points>
<intersection>-178 17</intersection>
<intersection>-137.5 1</intersection></vsegment>
<hsegment>
<ID>17</ID>
<points>-43,-178,-39.5,-178</points>
<connection>
<GID>161</GID>
<name>OUT_0</name></connection>
<intersection>-39.5 16</intersection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-41.5,-152,43.5,-152</points>
<connection>
<GID>45</GID>
<name>IN_1</name></connection>
<intersection>-41.5 15</intersection>
<intersection>24 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>24,-170.5,24,-152</points>
<intersection>-170.5 6</intersection>
<intersection>-164 4</intersection>
<intersection>-152 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>24,-164,37.5,-164</points>
<connection>
<GID>36</GID>
<name>IN_0</name></connection>
<intersection>24 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>24,-170.5,37.5,-170.5</points>
<connection>
<GID>37</GID>
<name>IN_0</name></connection>
<intersection>24 3</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>-41.5,-176,-41.5,-152</points>
<intersection>-176 16</intersection>
<intersection>-152 1</intersection></vsegment>
<hsegment>
<ID>16</ID>
<points>-43,-176,-41.5,-176</points>
<connection>
<GID>161</GID>
<name>OUT_1</name></connection>
<intersection>-41.5 15</intersection></hsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>43,-200.5,46,-200.5</points>
<connection>
<GID>65</GID>
<name>OUT</name></connection>
<connection>
<GID>66</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54,-199.5,54,-196</points>
<intersection>-199.5 2</intersection>
<intersection>-196 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>54,-196,57,-196</points>
<connection>
<GID>67</GID>
<name>IN_1</name></connection>
<intersection>54 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>52,-199.5,54,-199.5</points>
<connection>
<GID>66</GID>
<name>OUT</name></connection>
<intersection>54 0</intersection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>43,-194,57,-194</points>
<connection>
<GID>64</GID>
<name>OUT</name></connection>
<connection>
<GID>67</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>63,-195,66.5,-195</points>
<connection>
<GID>63</GID>
<name>N_in0</name></connection>
<intersection>63 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>63,-207.5,63,-195</points>
<connection>
<GID>67</GID>
<name>OUT</name></connection>
<intersection>-207.5 9</intersection>
<intersection>-195 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>42,-207.5,63,-207.5</points>
<connection>
<GID>83</GID>
<name>IN_0</name></connection>
<intersection>42 11</intersection>
<intersection>63 3</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>42,-227,42,-207.5</points>
<intersection>-227 12</intersection>
<intersection>-207.5 9</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>42,-227,45.5,-227</points>
<connection>
<GID>79</GID>
<name>IN_0</name></connection>
<intersection>42 11</intersection></hsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52,-184.5,52,-180</points>
<intersection>-184.5 1</intersection>
<intersection>-180 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>52,-184.5,55.5,-184.5</points>
<connection>
<GID>71</GID>
<name>IN_0</name></connection>
<intersection>52 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>49,-180,52,-180</points>
<connection>
<GID>70</GID>
<name>OUT</name></connection>
<intersection>52 0</intersection></hsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-25.5,-186.5,55.5,-186.5</points>
<connection>
<GID>71</GID>
<name>IN_1</name></connection>
<intersection>-25.5 8</intersection>
<intersection>35 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>35,-201.5,35,-186.5</points>
<intersection>-201.5 6</intersection>
<intersection>-195 4</intersection>
<intersection>-186.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>35,-195,37,-195</points>
<connection>
<GID>64</GID>
<name>IN_1</name></connection>
<intersection>35 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>35,-201.5,37,-201.5</points>
<connection>
<GID>65</GID>
<name>IN_1</name></connection>
<intersection>35 3</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>-25.5,-193,-25.5,-186.5</points>
<intersection>-193 9</intersection>
<intersection>-186.5 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>-43.5,-193,-25.5,-193</points>
<connection>
<GID>163</GID>
<name>OUT_2</name></connection>
<intersection>-25.5 8</intersection></hsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>61.5,-185.5,89,-185.5</points>
<connection>
<GID>71</GID>
<name>OUT</name></connection>
<connection>
<GID>72</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-33,-181,43,-181</points>
<connection>
<GID>70</GID>
<name>IN_1</name></connection>
<intersection>-33 15</intersection>
<intersection>36.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>36.5,-199.5,36.5,-181</points>
<intersection>-199.5 6</intersection>
<intersection>-193 4</intersection>
<intersection>-181 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>36.5,-193,37,-193</points>
<connection>
<GID>64</GID>
<name>IN_0</name></connection>
<intersection>36.5 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>36.5,-199.5,37,-199.5</points>
<connection>
<GID>65</GID>
<name>IN_0</name></connection>
<intersection>36.5 3</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>-33,-181,-33,-174</points>
<intersection>-181 1</intersection>
<intersection>-174 16</intersection></vsegment>
<hsegment>
<ID>16</ID>
<points>-43,-174,-33,-174</points>
<connection>
<GID>161</GID>
<name>OUT_2</name></connection>
<intersection>-33 15</intersection></hsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>42.5,-229,45.5,-229</points>
<connection>
<GID>78</GID>
<name>OUT</name></connection>
<connection>
<GID>79</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53.5,-228,53.5,-224.5</points>
<intersection>-228 2</intersection>
<intersection>-224.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>53.5,-224.5,56.5,-224.5</points>
<connection>
<GID>80</GID>
<name>IN_1</name></connection>
<intersection>53.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>51.5,-228,53.5,-228</points>
<connection>
<GID>79</GID>
<name>OUT</name></connection>
<intersection>53.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>42.5,-222.5,56.5,-222.5</points>
<connection>
<GID>77</GID>
<name>OUT</name></connection>
<connection>
<GID>80</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>47</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>51.5,-213,51.5,-208.5</points>
<intersection>-213 1</intersection>
<intersection>-208.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>51.5,-213,55,-213</points>
<connection>
<GID>84</GID>
<name>IN_0</name></connection>
<intersection>51.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>48.5,-208.5,51.5,-208.5</points>
<connection>
<GID>83</GID>
<name>OUT</name></connection>
<intersection>51.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-33,-215,55,-215</points>
<connection>
<GID>84</GID>
<name>IN_1</name></connection>
<intersection>-33 13</intersection>
<intersection>34.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>34.5,-230,34.5,-215</points>
<intersection>-230 6</intersection>
<intersection>-223.5 4</intersection>
<intersection>-215 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>34.5,-223.5,36.5,-223.5</points>
<connection>
<GID>77</GID>
<name>IN_1</name></connection>
<intersection>34.5 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>34.5,-230,36.5,-230</points>
<connection>
<GID>78</GID>
<name>IN_1</name></connection>
<intersection>34.5 3</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>-33,-215,-33,-191</points>
<intersection>-215 1</intersection>
<intersection>-191 14</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>-43.5,-191,-33,-191</points>
<connection>
<GID>163</GID>
<name>OUT_3</name></connection>
<intersection>-33 13</intersection></hsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>61,-214,89,-214</points>
<connection>
<GID>84</GID>
<name>OUT</name></connection>
<connection>
<GID>85</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-30.5,-209.5,42.5,-209.5</points>
<connection>
<GID>83</GID>
<name>IN_1</name></connection>
<intersection>-30.5 15</intersection>
<intersection>36 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>36,-228,36,-209.5</points>
<intersection>-228 6</intersection>
<intersection>-221.5 4</intersection>
<intersection>-209.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>36,-221.5,36.5,-221.5</points>
<connection>
<GID>77</GID>
<name>IN_0</name></connection>
<intersection>36 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>36,-228,36.5,-228</points>
<connection>
<GID>78</GID>
<name>IN_0</name></connection>
<intersection>36 3</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>-30.5,-209.5,-30.5,-172</points>
<intersection>-209.5 1</intersection>
<intersection>-172 16</intersection></vsegment>
<hsegment>
<ID>16</ID>
<points>-43,-172,-30.5,-172</points>
<connection>
<GID>161</GID>
<name>OUT_3</name></connection>
<intersection>-30.5 15</intersection></hsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<hsegment>
<ID>9</ID>
<points>42,-237.5,42.5,-237.5</points>
<connection>
<GID>96</GID>
<name>IN_0</name></connection>
<intersection>42 11</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>42,-257,42,-237.5</points>
<intersection>-257 12</intersection>
<intersection>-238 13</intersection>
<intersection>-237.5 9</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>42,-257,45.5,-257</points>
<connection>
<GID>92</GID>
<name>IN_0</name></connection>
<intersection>42 11</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>42,-238,65.5,-238</points>
<intersection>42 11</intersection>
<intersection>65.5 14</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>65.5,-238,65.5,-222.5</points>
<intersection>-238 13</intersection>
<intersection>-223.5 16</intersection>
<intersection>-222.5 15</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>65.5,-222.5,68.5,-222.5</points>
<connection>
<GID>76</GID>
<name>N_in0</name></connection>
<intersection>65.5 14</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>62.5,-223.5,65.5,-223.5</points>
<connection>
<GID>80</GID>
<name>OUT</name></connection>
<intersection>65.5 14</intersection></hsegment></shape></wire>
<wire>
<ID>52</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>42.5,-259,45.5,-259</points>
<connection>
<GID>91</GID>
<name>OUT</name></connection>
<connection>
<GID>92</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>53</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53.5,-258,53.5,-254.5</points>
<intersection>-258 2</intersection>
<intersection>-254.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>53.5,-254.5,56.5,-254.5</points>
<connection>
<GID>93</GID>
<name>IN_1</name></connection>
<intersection>53.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>51.5,-258,53.5,-258</points>
<connection>
<GID>92</GID>
<name>OUT</name></connection>
<intersection>53.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>54</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>42.5,-252.5,56.5,-252.5</points>
<connection>
<GID>90</GID>
<name>OUT</name></connection>
<connection>
<GID>93</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>56</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>51.5,-243,51.5,-238.5</points>
<intersection>-243 1</intersection>
<intersection>-238.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>51.5,-243,55,-243</points>
<connection>
<GID>97</GID>
<name>IN_0</name></connection>
<intersection>51.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>48.5,-238.5,51.5,-238.5</points>
<connection>
<GID>96</GID>
<name>OUT</name></connection>
<intersection>51.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>57</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-22,-245,55,-245</points>
<connection>
<GID>97</GID>
<name>IN_1</name></connection>
<intersection>-22 13</intersection>
<intersection>34.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>34.5,-260,34.5,-245</points>
<intersection>-260 6</intersection>
<intersection>-253.5 4</intersection>
<intersection>-245 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>34.5,-253.5,36.5,-253.5</points>
<connection>
<GID>90</GID>
<name>IN_1</name></connection>
<intersection>34.5 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>34.5,-260,36.5,-260</points>
<connection>
<GID>91</GID>
<name>IN_1</name></connection>
<intersection>34.5 3</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>-22,-299.5,-22,-245</points>
<intersection>-299.5 14</intersection>
<intersection>-245 1</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>-48.5,-299.5,-22,-299.5</points>
<connection>
<GID>167</GID>
<name>OUT_0</name></connection>
<intersection>-22 13</intersection></hsegment></shape></wire>
<wire>
<ID>58</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>61,-244,88.5,-244</points>
<connection>
<GID>97</GID>
<name>OUT</name></connection>
<connection>
<GID>98</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>59</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-33,-239.5,42.5,-239.5</points>
<connection>
<GID>96</GID>
<name>IN_1</name></connection>
<intersection>-33 13</intersection>
<intersection>36 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>36,-258,36,-239.5</points>
<intersection>-258 6</intersection>
<intersection>-251.5 4</intersection>
<intersection>-239.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>36,-251.5,36.5,-251.5</points>
<connection>
<GID>90</GID>
<name>IN_0</name></connection>
<intersection>36 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>36,-258,36.5,-258</points>
<connection>
<GID>91</GID>
<name>IN_0</name></connection>
<intersection>36 3</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>-33,-281.5,-33,-239.5</points>
<intersection>-281.5 14</intersection>
<intersection>-239.5 1</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>-48,-281.5,-33,-281.5</points>
<connection>
<GID>165</GID>
<name>OUT_0</name></connection>
<intersection>-33 13</intersection></hsegment></shape></wire>
<wire>
<ID>60</ID>
<shape>
<hsegment>
<ID>9</ID>
<points>38.5,-266.5,65.5,-266.5</points>
<connection>
<GID>109</GID>
<name>IN_0</name></connection>
<intersection>38.5 11</intersection>
<intersection>65.5 14</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>38.5,-286,38.5,-266.5</points>
<intersection>-286 12</intersection>
<intersection>-266.5 9</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>38.5,-286,42,-286</points>
<connection>
<GID>105</GID>
<name>IN_0</name></connection>
<intersection>38.5 11</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>65.5,-266.5,65.5,-252.5</points>
<intersection>-266.5 9</intersection>
<intersection>-253.5 16</intersection>
<intersection>-252.5 15</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>65.5,-252.5,68.5,-252.5</points>
<connection>
<GID>89</GID>
<name>N_in0</name></connection>
<intersection>65.5 14</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>62.5,-253.5,65.5,-253.5</points>
<connection>
<GID>93</GID>
<name>OUT</name></connection>
<intersection>65.5 14</intersection></hsegment></shape></wire>
<wire>
<ID>61</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>39,-288,42,-288</points>
<connection>
<GID>104</GID>
<name>OUT</name></connection>
<connection>
<GID>105</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>62</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50,-287,50,-283.5</points>
<intersection>-287 2</intersection>
<intersection>-283.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50,-283.5,53,-283.5</points>
<connection>
<GID>106</GID>
<name>IN_1</name></connection>
<intersection>50 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>48,-287,50,-287</points>
<connection>
<GID>105</GID>
<name>OUT</name></connection>
<intersection>50 0</intersection></hsegment></shape></wire>
<wire>
<ID>63</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>39,-281.5,53,-281.5</points>
<connection>
<GID>103</GID>
<name>OUT</name></connection>
<connection>
<GID>106</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>48,-272,48,-267.5</points>
<intersection>-272 1</intersection>
<intersection>-267.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>48,-272,51.5,-272</points>
<connection>
<GID>110</GID>
<name>IN_0</name></connection>
<intersection>48 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>45,-267.5,48,-267.5</points>
<connection>
<GID>109</GID>
<name>OUT</name></connection>
<intersection>48 0</intersection></hsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-27,-274,51.5,-274</points>
<connection>
<GID>110</GID>
<name>IN_1</name></connection>
<intersection>-27 17</intersection>
<intersection>31 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>31,-289,31,-274</points>
<intersection>-289 6</intersection>
<intersection>-282.5 4</intersection>
<intersection>-274 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>31,-282.5,33,-282.5</points>
<connection>
<GID>103</GID>
<name>IN_1</name></connection>
<intersection>31 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>31,-289,33,-289</points>
<connection>
<GID>104</GID>
<name>IN_1</name></connection>
<intersection>31 3</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>-27,-297.5,-27,-274</points>
<intersection>-297.5 18</intersection>
<intersection>-274 1</intersection></vsegment>
<hsegment>
<ID>18</ID>
<points>-48.5,-297.5,-27,-297.5</points>
<connection>
<GID>167</GID>
<name>OUT_1</name></connection>
<intersection>-27 17</intersection></hsegment></shape></wire>
<wire>
<ID>67</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>57.5,-273,89,-273</points>
<connection>
<GID>110</GID>
<name>OUT</name></connection>
<connection>
<GID>111</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>68</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-38,-268.5,39,-268.5</points>
<connection>
<GID>109</GID>
<name>IN_1</name></connection>
<intersection>-38 14</intersection>
<intersection>32.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>32.5,-287,32.5,-268.5</points>
<intersection>-287 6</intersection>
<intersection>-280.5 4</intersection>
<intersection>-268.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>32.5,-280.5,33,-280.5</points>
<connection>
<GID>103</GID>
<name>IN_0</name></connection>
<intersection>32.5 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>32.5,-287,33,-287</points>
<connection>
<GID>104</GID>
<name>IN_0</name></connection>
<intersection>32.5 3</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>-38,-279.5,-38,-268.5</points>
<intersection>-279.5 15</intersection>
<intersection>-268.5 1</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>-48,-279.5,-38,-279.5</points>
<connection>
<GID>165</GID>
<name>OUT_1</name></connection>
<intersection>-38 14</intersection></hsegment></shape></wire>
<wire>
<ID>69</ID>
<shape>
<hsegment>
<ID>9</ID>
<points>36.5,-295,59,-295</points>
<connection>
<GID>122</GID>
<name>IN_0</name></connection>
<intersection>36.5 11</intersection>
<intersection>59 13</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>36.5,-314.5,36.5,-295</points>
<intersection>-314.5 12</intersection>
<intersection>-295 9</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>36.5,-314.5,40,-314.5</points>
<connection>
<GID>118</GID>
<name>IN_0</name></connection>
<intersection>36.5 11</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>59,-295,59,-282.5</points>
<connection>
<GID>106</GID>
<name>OUT</name></connection>
<intersection>-295 9</intersection>
<intersection>-282.5 15</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>59,-282.5,66,-282.5</points>
<connection>
<GID>102</GID>
<name>N_in0</name></connection>
<intersection>59 13</intersection></hsegment></shape></wire>
<wire>
<ID>70</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>37,-316.5,40,-316.5</points>
<connection>
<GID>117</GID>
<name>OUT</name></connection>
<connection>
<GID>118</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>71</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>48,-315.5,48,-312</points>
<intersection>-315.5 2</intersection>
<intersection>-312 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>48,-312,51,-312</points>
<connection>
<GID>119</GID>
<name>IN_1</name></connection>
<intersection>48 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>46,-315.5,48,-315.5</points>
<connection>
<GID>118</GID>
<name>OUT</name></connection>
<intersection>48 0</intersection></hsegment></shape></wire>
<wire>
<ID>72</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>37,-310,51,-310</points>
<connection>
<GID>116</GID>
<name>OUT</name></connection>
<connection>
<GID>119</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>74</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>46,-300.5,46,-296</points>
<intersection>-300.5 1</intersection>
<intersection>-296 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>46,-300.5,49.5,-300.5</points>
<connection>
<GID>123</GID>
<name>IN_0</name></connection>
<intersection>46 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>43,-296,46,-296</points>
<connection>
<GID>122</GID>
<name>OUT</name></connection>
<intersection>46 0</intersection></hsegment></shape></wire>
<wire>
<ID>75</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-43,-302.5,49.5,-302.5</points>
<connection>
<GID>123</GID>
<name>IN_1</name></connection>
<intersection>-43 18</intersection>
<intersection>29 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>29,-317.5,29,-302.5</points>
<intersection>-317.5 6</intersection>
<intersection>-311 4</intersection>
<intersection>-302.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>29,-311,31,-311</points>
<connection>
<GID>116</GID>
<name>IN_1</name></connection>
<intersection>29 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>29,-317.5,31,-317.5</points>
<connection>
<GID>117</GID>
<name>IN_1</name></connection>
<intersection>29 3</intersection></hsegment>
<vsegment>
<ID>18</ID>
<points>-43,-302.5,-43,-295.5</points>
<intersection>-302.5 1</intersection>
<intersection>-295.5 19</intersection></vsegment>
<hsegment>
<ID>19</ID>
<points>-48.5,-295.5,-43,-295.5</points>
<connection>
<GID>167</GID>
<name>OUT_2</name></connection>
<intersection>-43 18</intersection></hsegment></shape></wire>
<wire>
<ID>76</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>55.5,-301.5,89,-301.5</points>
<connection>
<GID>123</GID>
<name>OUT</name></connection>
<connection>
<GID>124</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>77</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-40.5,-297,37,-297</points>
<connection>
<GID>122</GID>
<name>IN_1</name></connection>
<intersection>-40.5 14</intersection>
<intersection>30.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>30.5,-315.5,30.5,-297</points>
<intersection>-315.5 6</intersection>
<intersection>-309 4</intersection>
<intersection>-297 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>30.5,-309,31,-309</points>
<connection>
<GID>116</GID>
<name>IN_0</name></connection>
<intersection>30.5 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>30.5,-315.5,31,-315.5</points>
<connection>
<GID>117</GID>
<name>IN_0</name></connection>
<intersection>30.5 3</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>-40.5,-297,-40.5,-277.5</points>
<intersection>-297 1</intersection>
<intersection>-277.5 15</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>-48,-277.5,-40.5,-277.5</points>
<connection>
<GID>165</GID>
<name>OUT_2</name></connection>
<intersection>-40.5 14</intersection></hsegment></shape></wire>
<wire>
<ID>78</ID>
<shape>
<hsegment>
<ID>9</ID>
<points>36,-324,56.5,-324</points>
<connection>
<GID>135</GID>
<name>IN_0</name></connection>
<intersection>36 11</intersection>
<intersection>56.5 13</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>36,-343.5,36,-324</points>
<intersection>-343.5 12</intersection>
<intersection>-324 9</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>36,-343.5,39.5,-343.5</points>
<connection>
<GID>131</GID>
<name>IN_0</name></connection>
<intersection>36 11</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>56.5,-324,56.5,-311</points>
<intersection>-324 9</intersection>
<intersection>-311 15</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>56.5,-311,63,-311</points>
<connection>
<GID>119</GID>
<name>OUT</name></connection>
<connection>
<GID>115</GID>
<name>N_in0</name></connection>
<intersection>56.5 13</intersection></hsegment></shape></wire>
<wire>
<ID>79</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>36.5,-345.5,39.5,-345.5</points>
<connection>
<GID>130</GID>
<name>OUT</name></connection>
<connection>
<GID>131</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>80</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47.5,-344.5,47.5,-341</points>
<intersection>-344.5 2</intersection>
<intersection>-341 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47.5,-341,50.5,-341</points>
<connection>
<GID>132</GID>
<name>IN_1</name></connection>
<intersection>47.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>45.5,-344.5,47.5,-344.5</points>
<connection>
<GID>131</GID>
<name>OUT</name></connection>
<intersection>47.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>81</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>36.5,-339,50.5,-339</points>
<connection>
<GID>129</GID>
<name>OUT</name></connection>
<connection>
<GID>132</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>83</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45.5,-329.5,45.5,-325</points>
<intersection>-329.5 1</intersection>
<intersection>-325 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>45.5,-329.5,49,-329.5</points>
<connection>
<GID>136</GID>
<name>IN_0</name></connection>
<intersection>45.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>42.5,-325,45.5,-325</points>
<connection>
<GID>135</GID>
<name>OUT</name></connection>
<intersection>45.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>84</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-35.5,-331.5,49,-331.5</points>
<connection>
<GID>136</GID>
<name>IN_1</name></connection>
<intersection>-35.5 16</intersection>
<intersection>28.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>28.5,-346.5,28.5,-331.5</points>
<intersection>-346.5 6</intersection>
<intersection>-340 4</intersection>
<intersection>-331.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>28.5,-340,30.5,-340</points>
<connection>
<GID>129</GID>
<name>IN_1</name></connection>
<intersection>28.5 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>28.5,-346.5,30.5,-346.5</points>
<connection>
<GID>130</GID>
<name>IN_1</name></connection>
<intersection>28.5 3</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>-35.5,-331.5,-35.5,-293.5</points>
<intersection>-331.5 1</intersection>
<intersection>-293.5 17</intersection></vsegment>
<hsegment>
<ID>17</ID>
<points>-48.5,-293.5,-35.5,-293.5</points>
<connection>
<GID>167</GID>
<name>OUT_3</name></connection>
<intersection>-35.5 16</intersection></hsegment></shape></wire>
<wire>
<ID>85</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>55,-330.5,88.5,-330.5</points>
<connection>
<GID>136</GID>
<name>OUT</name></connection>
<connection>
<GID>137</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>86</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-25,-326,36.5,-326</points>
<connection>
<GID>135</GID>
<name>IN_1</name></connection>
<intersection>-25 14</intersection>
<intersection>30 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>30,-344.5,30,-326</points>
<intersection>-344.5 6</intersection>
<intersection>-338 4</intersection>
<intersection>-326 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>30,-338,30.5,-338</points>
<connection>
<GID>129</GID>
<name>IN_0</name></connection>
<intersection>30 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>30,-344.5,30.5,-344.5</points>
<connection>
<GID>130</GID>
<name>IN_0</name></connection>
<intersection>30 3</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>-25,-326,-25,-275.5</points>
<intersection>-326 1</intersection>
<intersection>-275.5 15</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>-48,-275.5,-25,-275.5</points>
<connection>
<GID>165</GID>
<name>OUT_3</name></connection>
<intersection>-25 14</intersection></hsegment></shape></wire>
<wire>
<ID>87</ID>
<shape>
<hsegment>
<ID>15</ID>
<points>56.5,-340,77.5,-340</points>
<connection>
<GID>132</GID>
<name>OUT</name></connection>
<connection>
<GID>128</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>96</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>67.5,-167,67.5,-166</points>
<connection>
<GID>35</GID>
<name>N_in2</name></connection>
<intersection>-166 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>67.5,-166,68.5,-166</points>
<connection>
<GID>35</GID>
<name>N_in1</name></connection>
<intersection>67.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>99</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>79.5,-340,169.5,-340</points>
<connection>
<GID>128</GID>
<name>N_in1</name></connection>
<connection>
<GID>171</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>100</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>137,-229,137,-138.5</points>
<intersection>-229 1</intersection>
<intersection>-138.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>137,-229,176,-229</points>
<connection>
<GID>169</GID>
<name>IN_0</name></connection>
<intersection>137 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>90,-138.5,137,-138.5</points>
<connection>
<GID>11</GID>
<name>N_in1</name></connection>
<intersection>137 0</intersection></hsegment></shape></wire>
<wire>
<ID>101</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>133.5,-228,133.5,-156.5</points>
<intersection>-228 1</intersection>
<intersection>-156.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>133.5,-228,176,-228</points>
<connection>
<GID>169</GID>
<name>IN_1</name></connection>
<intersection>133.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>90.5,-156.5,133.5,-156.5</points>
<connection>
<GID>48</GID>
<name>N_in1</name></connection>
<intersection>133.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>102</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>129.5,-227,129.5,-185.5</points>
<intersection>-227 1</intersection>
<intersection>-185.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>129.5,-227,176,-227</points>
<connection>
<GID>169</GID>
<name>IN_2</name></connection>
<intersection>129.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>91,-185.5,129.5,-185.5</points>
<connection>
<GID>72</GID>
<name>N_in1</name></connection>
<intersection>129.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>103</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>127,-226,127,-214</points>
<intersection>-226 1</intersection>
<intersection>-214 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>127,-226,176,-226</points>
<connection>
<GID>169</GID>
<name>IN_3</name></connection>
<intersection>127 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>91,-214,127,-214</points>
<connection>
<GID>85</GID>
<name>N_in1</name></connection>
<intersection>127 0</intersection></hsegment></shape></wire>
<wire>
<ID>104</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>125,-244,125,-225</points>
<intersection>-244 2</intersection>
<intersection>-225 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>125,-225,176,-225</points>
<connection>
<GID>169</GID>
<name>IN_4</name></connection>
<intersection>125 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>90.5,-244,125,-244</points>
<connection>
<GID>98</GID>
<name>N_in1</name></connection>
<intersection>125 0</intersection></hsegment></shape></wire>
<wire>
<ID>105</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>121,-273,121,-224</points>
<intersection>-273 2</intersection>
<intersection>-224 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>121,-224,176,-224</points>
<connection>
<GID>169</GID>
<name>IN_5</name></connection>
<intersection>121 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>91,-273,121,-273</points>
<connection>
<GID>111</GID>
<name>N_in1</name></connection>
<intersection>121 0</intersection></hsegment></shape></wire>
<wire>
<ID>106</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>116,-301.5,116,-223</points>
<intersection>-301.5 2</intersection>
<intersection>-223 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>116,-223,176,-223</points>
<connection>
<GID>169</GID>
<name>IN_6</name></connection>
<intersection>116 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>91,-301.5,116,-301.5</points>
<connection>
<GID>124</GID>
<name>N_in1</name></connection>
<intersection>116 0</intersection></hsegment></shape></wire>
<wire>
<ID>107</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>110,-330.5,110,-222</points>
<intersection>-330.5 2</intersection>
<intersection>-222 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>110,-222,176,-222</points>
<connection>
<GID>169</GID>
<name>IN_7</name></connection>
<intersection>110 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>90.5,-330.5,110,-330.5</points>
<connection>
<GID>137</GID>
<name>N_in1</name></connection>
<intersection>110 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,4.04748e-006,177.8,-91.7</PageViewport></page 1>
<page 2>
<PageViewport>0,4.04748e-006,177.8,-91.7</PageViewport></page 2>
<page 3>
<PageViewport>0,4.04748e-006,177.8,-91.7</PageViewport></page 3>
<page 4>
<PageViewport>0,4.04748e-006,177.8,-91.7</PageViewport></page 4>
<page 5>
<PageViewport>0,4.04748e-006,177.8,-91.7</PageViewport></page 5>
<page 6>
<PageViewport>0,4.04748e-006,177.8,-91.7</PageViewport></page 6>
<page 7>
<PageViewport>0,4.04748e-006,177.8,-91.7</PageViewport></page 7>
<page 8>
<PageViewport>0,4.04748e-006,177.8,-91.7</PageViewport></page 8>
<page 9>
<PageViewport>0,4.04748e-006,177.8,-91.7</PageViewport></page 9></circuit>