<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-10.8311,-76.6697,170.471,-170.176</PageViewport>
<gate>
<ID>2</ID>
<type>AA_LABEL</type>
<position>65,-85</position>
<gparam>LABEL_TEXT 4bit Encoder</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>8</ID>
<type>AA_TOGGLE</type>
<position>46.5,-95.5</position>
<output>
<ID>OUT_0</ID>59 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>10</ID>
<type>AA_TOGGLE</type>
<position>46.5,-98.5</position>
<output>
<ID>OUT_0</ID>52 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>12</ID>
<type>AA_TOGGLE</type>
<position>46.5,-102</position>
<output>
<ID>OUT_0</ID>50 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>14</ID>
<type>AA_TOGGLE</type>
<position>46.5,-106</position>
<output>
<ID>OUT_0</ID>51 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>17</ID>
<type>AA_LABEL</type>
<position>42,-94</position>
<gparam>LABEL_TEXT D0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>18</ID>
<type>AA_LABEL</type>
<position>42,-98</position>
<gparam>LABEL_TEXT D1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>19</ID>
<type>AA_LABEL</type>
<position>42,-102</position>
<gparam>LABEL_TEXT D2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>20</ID>
<type>AA_LABEL</type>
<position>42,-105.5</position>
<gparam>LABEL_TEXT D3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>34</ID>
<type>AA_TOGGLE</type>
<position>38,-127</position>
<output>
<ID>OUT_0</ID>65 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>35</ID>
<type>AA_TOGGLE</type>
<position>38.5,-131.5</position>
<output>
<ID>OUT_0</ID>67 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>36</ID>
<type>AA_TOGGLE</type>
<position>38.5,-135.5</position>
<output>
<ID>OUT_0</ID>86 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>37</ID>
<type>AA_TOGGLE</type>
<position>38.5,-139.5</position>
<output>
<ID>OUT_0</ID>74 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>38</ID>
<type>AA_LABEL</type>
<position>34,-127</position>
<gparam>LABEL_TEXT I0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>39</ID>
<type>AA_LABEL</type>
<position>34,-131</position>
<gparam>LABEL_TEXT I1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>40</ID>
<type>AA_LABEL</type>
<position>34,-135</position>
<gparam>LABEL_TEXT I2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>41</ID>
<type>AA_LABEL</type>
<position>34,-138.5</position>
<gparam>LABEL_TEXT I3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>48</ID>
<type>AA_TOGGLE</type>
<position>38.5,-144</position>
<output>
<ID>OUT_0</ID>83 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>49</ID>
<type>AA_TOGGLE</type>
<position>38.5,-149</position>
<output>
<ID>OUT_0</ID>69 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>50</ID>
<type>AA_TOGGLE</type>
<position>38.5,-153</position>
<output>
<ID>OUT_0</ID>76 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>51</ID>
<type>AA_TOGGLE</type>
<position>38.5,-157</position>
<output>
<ID>OUT_0</ID>70 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>52</ID>
<type>AA_LABEL</type>
<position>34,-144.5</position>
<gparam>LABEL_TEXT I4</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>53</ID>
<type>AA_LABEL</type>
<position>34,-148.5</position>
<gparam>LABEL_TEXT I5</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>54</ID>
<type>AA_LABEL</type>
<position>34,-152.5</position>
<gparam>LABEL_TEXT I6</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>55</ID>
<type>AA_LABEL</type>
<position>34,-156</position>
<gparam>LABEL_TEXT I7</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>61</ID>
<type>AA_LABEL</type>
<position>111,-129.5</position>
<gparam>LABEL_TEXT X</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>62</ID>
<type>GA_LED</type>
<position>111,-132.5</position>
<input>
<ID>N_in0</ID>79 </input>
<input>
<ID>N_in2</ID>93 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>63</ID>
<type>AA_LABEL</type>
<position>108,-140.5</position>
<gparam>LABEL_TEXT y</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>64</ID>
<type>GA_LED</type>
<position>108.5,-144</position>
<input>
<ID>N_in0</ID>80 </input>
<input>
<ID>N_in3</ID>92 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>65</ID>
<type>AA_LABEL</type>
<position>103,-150.5</position>
<gparam>LABEL_TEXT z</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>66</ID>
<type>GA_LED</type>
<position>103.5,-154</position>
<input>
<ID>N_in0</ID>81 </input>
<input>
<ID>N_in1</ID>91 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>98</ID>
<type>AE_OR2</type>
<position>65,-97</position>
<input>
<ID>IN_0</ID>50 </input>
<input>
<ID>IN_1</ID>51 </input>
<output>
<ID>OUT</ID>61 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>100</ID>
<type>AE_OR2</type>
<position>65.5,-104.5</position>
<input>
<ID>IN_0</ID>52 </input>
<input>
<ID>IN_1</ID>51 </input>
<output>
<ID>OUT</ID>62 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>110</ID>
<type>AA_AND2</type>
<position>75.5,-98</position>
<input>
<ID>IN_0</ID>60 </input>
<input>
<ID>IN_1</ID>61 </input>
<output>
<ID>OUT</ID>63 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>112</ID>
<type>AA_AND2</type>
<position>76,-104.5</position>
<input>
<ID>IN_0</ID>62 </input>
<input>
<ID>IN_1</ID>60 </input>
<output>
<ID>OUT</ID>64 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>114</ID>
<type>AA_INVERTER</type>
<position>67,-91</position>
<input>
<ID>IN_0</ID>59 </input>
<output>
<ID>OUT_0</ID>60 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>115</ID>
<type>AA_LABEL</type>
<position>87.5,-94</position>
<gparam>LABEL_TEXT X</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>116</ID>
<type>GA_LED</type>
<position>88,-97.5</position>
<input>
<ID>N_in0</ID>63 </input>
<input>
<ID>N_in1</ID>97 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>117</ID>
<type>AA_LABEL</type>
<position>87.5,-101</position>
<gparam>LABEL_TEXT y</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>118</ID>
<type>GA_LED</type>
<position>88,-104.5</position>
<input>
<ID>N_in0</ID>64 </input>
<input>
<ID>N_in1</ID>96 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>120</ID>
<type>AE_OR2</type>
<position>61,-129.5</position>
<input>
<ID>IN_0</ID>67 </input>
<input>
<ID>IN_1</ID>74 </input>
<output>
<ID>OUT</ID>71 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>122</ID>
<type>AE_OR2</type>
<position>70.5,-130.5</position>
<input>
<ID>IN_0</ID>71 </input>
<input>
<ID>IN_1</ID>69 </input>
<output>
<ID>OUT</ID>72 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>124</ID>
<type>AE_OR2</type>
<position>81,-131.5</position>
<input>
<ID>IN_0</ID>72 </input>
<input>
<ID>IN_1</ID>70 </input>
<output>
<ID>OUT</ID>73 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>126</ID>
<type>AA_AND2</type>
<position>92.5,-132.5</position>
<input>
<ID>IN_0</ID>73 </input>
<input>
<ID>IN_1</ID>66 </input>
<output>
<ID>OUT</ID>79 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>127</ID>
<type>AA_INVERTER</type>
<position>73.5,-123.5</position>
<input>
<ID>IN_0</ID>65 </input>
<output>
<ID>OUT_0</ID>66 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>128</ID>
<type>AE_OR2</type>
<position>61.5,-141</position>
<input>
<ID>IN_0</ID>86 </input>
<input>
<ID>IN_1</ID>74 </input>
<output>
<ID>OUT</ID>75 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>129</ID>
<type>AE_OR2</type>
<position>70.5,-142</position>
<input>
<ID>IN_0</ID>75 </input>
<input>
<ID>IN_1</ID>76 </input>
<output>
<ID>OUT</ID>77 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>130</ID>
<type>AE_OR2</type>
<position>80.5,-143</position>
<input>
<ID>IN_0</ID>77 </input>
<input>
<ID>IN_1</ID>70 </input>
<output>
<ID>OUT</ID>78 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>131</ID>
<type>AA_AND2</type>
<position>93,-144</position>
<input>
<ID>IN_0</ID>78 </input>
<input>
<ID>IN_1</ID>66 </input>
<output>
<ID>OUT</ID>80 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>132</ID>
<type>AE_OR2</type>
<position>61.5,-151</position>
<input>
<ID>IN_0</ID>83 </input>
<input>
<ID>IN_1</ID>69 </input>
<output>
<ID>OUT</ID>84 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>133</ID>
<type>AE_OR2</type>
<position>70.5,-152</position>
<input>
<ID>IN_0</ID>84 </input>
<input>
<ID>IN_1</ID>76 </input>
<output>
<ID>OUT</ID>85 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>134</ID>
<type>AE_OR2</type>
<position>81,-153</position>
<input>
<ID>IN_0</ID>85 </input>
<input>
<ID>IN_1</ID>70 </input>
<output>
<ID>OUT</ID>82 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>135</ID>
<type>AA_AND2</type>
<position>93,-154</position>
<input>
<ID>IN_0</ID>82 </input>
<input>
<ID>IN_1</ID>66 </input>
<output>
<ID>OUT</ID>81 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>139</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>121,-140</position>
<input>
<ID>IN_0</ID>93 </input>
<input>
<ID>IN_1</ID>92 </input>
<input>
<ID>IN_2</ID>91 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>142</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>100.5,-100</position>
<input>
<ID>IN_0</ID>96 </input>
<input>
<ID>IN_1</ID>97 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>143</ID>
<type>AA_LABEL</type>
<position>63.5,-118.5</position>
<gparam>LABEL_TEXT 8bit Encoder</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>50</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>55,-102,55,-96</points>
<intersection>-102 2</intersection>
<intersection>-96 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>55,-96,62,-96</points>
<connection>
<GID>98</GID>
<name>IN_0</name></connection>
<intersection>55 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>48.5,-102,55,-102</points>
<connection>
<GID>12</GID>
<name>OUT_0</name></connection>
<intersection>55 0</intersection></hsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56.5,-106,56.5,-98</points>
<intersection>-106 2</intersection>
<intersection>-98 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>56.5,-98,62,-98</points>
<connection>
<GID>98</GID>
<name>IN_1</name></connection>
<intersection>56.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>48.5,-106,62.5,-106</points>
<connection>
<GID>14</GID>
<name>OUT_0</name></connection>
<intersection>56.5 0</intersection>
<intersection>62.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>62.5,-106,62.5,-105.5</points>
<connection>
<GID>100</GID>
<name>IN_1</name></connection>
<intersection>-106 2</intersection></vsegment></shape></wire>
<wire>
<ID>52</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>55.5,-103.5,55.5,-98.5</points>
<intersection>-103.5 1</intersection>
<intersection>-98.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>55.5,-103.5,62.5,-103.5</points>
<connection>
<GID>100</GID>
<name>IN_0</name></connection>
<intersection>55.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>48.5,-98.5,55.5,-98.5</points>
<connection>
<GID>10</GID>
<name>OUT_0</name></connection>
<intersection>55.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>59</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56,-95.5,56,-91</points>
<intersection>-95.5 2</intersection>
<intersection>-91 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>56,-91,64,-91</points>
<connection>
<GID>114</GID>
<name>IN_0</name></connection>
<intersection>56 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>48.5,-95.5,56,-95.5</points>
<connection>
<GID>8</GID>
<name>OUT_0</name></connection>
<intersection>56 0</intersection></hsegment></shape></wire>
<wire>
<ID>60</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>71,-97,71,-91</points>
<intersection>-97 1</intersection>
<intersection>-91 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>71,-97,72.5,-97</points>
<connection>
<GID>110</GID>
<name>IN_0</name></connection>
<intersection>71 0</intersection>
<intersection>71.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>70,-91,71,-91</points>
<connection>
<GID>114</GID>
<name>OUT_0</name></connection>
<intersection>71 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>71.5,-105.5,71.5,-97</points>
<intersection>-105.5 4</intersection>
<intersection>-97 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>71.5,-105.5,73,-105.5</points>
<connection>
<GID>112</GID>
<name>IN_1</name></connection>
<intersection>71.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>61</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>70,-99,70,-97</points>
<intersection>-99 1</intersection>
<intersection>-97 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>70,-99,72.5,-99</points>
<connection>
<GID>110</GID>
<name>IN_1</name></connection>
<intersection>70 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>68,-97,70,-97</points>
<connection>
<GID>98</GID>
<name>OUT</name></connection>
<intersection>70 0</intersection></hsegment></shape></wire>
<wire>
<ID>62</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>70.5,-104.5,70.5,-103.5</points>
<intersection>-104.5 2</intersection>
<intersection>-103.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>70.5,-103.5,73,-103.5</points>
<connection>
<GID>112</GID>
<name>IN_0</name></connection>
<intersection>70.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>68.5,-104.5,70.5,-104.5</points>
<connection>
<GID>100</GID>
<name>OUT</name></connection>
<intersection>70.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>63</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>82.5,-98,82.5,-97.5</points>
<intersection>-98 2</intersection>
<intersection>-97.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>82.5,-97.5,87,-97.5</points>
<connection>
<GID>116</GID>
<name>N_in0</name></connection>
<intersection>82.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>78.5,-98,82.5,-98</points>
<connection>
<GID>110</GID>
<name>OUT</name></connection>
<intersection>82.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>64</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>79,-104.5,87,-104.5</points>
<connection>
<GID>112</GID>
<name>OUT</name></connection>
<connection>
<GID>118</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>55.5,-127,55.5,-123.5</points>
<intersection>-127 2</intersection>
<intersection>-123.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>55.5,-123.5,70.5,-123.5</points>
<connection>
<GID>127</GID>
<name>IN_0</name></connection>
<intersection>55.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>40,-127,55.5,-127</points>
<connection>
<GID>34</GID>
<name>OUT_0</name></connection>
<intersection>55.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>86,-133.5,86,-123.5</points>
<intersection>-133.5 1</intersection>
<intersection>-123.5 7</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>86,-133.5,89.5,-133.5</points>
<connection>
<GID>126</GID>
<name>IN_1</name></connection>
<intersection>86 0</intersection>
<intersection>87.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>87.5,-155,87.5,-133.5</points>
<intersection>-155 5</intersection>
<intersection>-145 6</intersection>
<intersection>-133.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>87.5,-155,90,-155</points>
<connection>
<GID>135</GID>
<name>IN_1</name></connection>
<intersection>87.5 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>87.5,-145,90,-145</points>
<connection>
<GID>131</GID>
<name>IN_1</name></connection>
<intersection>87.5 3</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>76.5,-123.5,86,-123.5</points>
<connection>
<GID>127</GID>
<name>OUT_0</name></connection>
<intersection>86 0</intersection></hsegment></shape></wire>
<wire>
<ID>67</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49,-131.5,49,-128.5</points>
<intersection>-131.5 2</intersection>
<intersection>-128.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>49,-128.5,58,-128.5</points>
<connection>
<GID>120</GID>
<name>IN_0</name></connection>
<intersection>49 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>40.5,-131.5,49,-131.5</points>
<connection>
<GID>35</GID>
<name>OUT_0</name></connection>
<intersection>49 0</intersection></hsegment></shape></wire>
<wire>
<ID>69</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54,-152,54,-131.5</points>
<intersection>-152 3</intersection>
<intersection>-149 2</intersection>
<intersection>-131.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>54,-131.5,67.5,-131.5</points>
<connection>
<GID>122</GID>
<name>IN_1</name></connection>
<intersection>54 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>40.5,-149,54,-149</points>
<connection>
<GID>49</GID>
<name>OUT_0</name></connection>
<intersection>54 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>54,-152,58.5,-152</points>
<connection>
<GID>132</GID>
<name>IN_1</name></connection>
<intersection>54 0</intersection></hsegment></shape></wire>
<wire>
<ID>70</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>55.5,-157,55.5,-132.5</points>
<intersection>-157 2</intersection>
<intersection>-132.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>55.5,-132.5,78,-132.5</points>
<connection>
<GID>124</GID>
<name>IN_1</name></connection>
<intersection>55.5 0</intersection>
<intersection>76.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>40.5,-157,55.5,-157</points>
<connection>
<GID>51</GID>
<name>OUT_0</name></connection>
<intersection>55.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>76.5,-144,76.5,-132.5</points>
<intersection>-144 4</intersection>
<intersection>-132.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>76.5,-144,77.5,-144</points>
<connection>
<GID>130</GID>
<name>IN_1</name></connection>
<intersection>76.5 3</intersection>
<intersection>77 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>77,-154,77,-144</points>
<intersection>-154 6</intersection>
<intersection>-144 4</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>77,-154,78,-154</points>
<connection>
<GID>134</GID>
<name>IN_1</name></connection>
<intersection>77 5</intersection></hsegment></shape></wire>
<wire>
<ID>71</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>64,-129.5,67.5,-129.5</points>
<connection>
<GID>120</GID>
<name>OUT</name></connection>
<connection>
<GID>122</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>72</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73.5,-130.5,78,-130.5</points>
<connection>
<GID>122</GID>
<name>OUT</name></connection>
<connection>
<GID>124</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>73</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>84,-131.5,89.5,-131.5</points>
<connection>
<GID>124</GID>
<name>OUT</name></connection>
<connection>
<GID>126</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>74</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49.5,-142,49.5,-139.5</points>
<intersection>-142 2</intersection>
<intersection>-139.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>40.5,-139.5,49.5,-139.5</points>
<connection>
<GID>37</GID>
<name>OUT_0</name></connection>
<intersection>49.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>49.5,-142,58.5,-142</points>
<connection>
<GID>128</GID>
<name>IN_1</name></connection>
<intersection>49.5 0</intersection>
<intersection>57 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>57,-142,57,-130.5</points>
<intersection>-142 2</intersection>
<intersection>-130.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>57,-130.5,58,-130.5</points>
<connection>
<GID>120</GID>
<name>IN_1</name></connection>
<intersection>57 3</intersection></hsegment></shape></wire>
<wire>
<ID>75</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>64.5,-141,67.5,-141</points>
<connection>
<GID>128</GID>
<name>OUT</name></connection>
<connection>
<GID>129</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>76</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52.5,-153,52.5,-143</points>
<intersection>-153 1</intersection>
<intersection>-143 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>40.5,-153,52.5,-153</points>
<connection>
<GID>50</GID>
<name>OUT_0</name></connection>
<intersection>52.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>52.5,-143,67.5,-143</points>
<connection>
<GID>129</GID>
<name>IN_1</name></connection>
<intersection>52.5 0</intersection>
<intersection>65.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>65.5,-153,65.5,-143</points>
<intersection>-153 4</intersection>
<intersection>-143 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>65.5,-153,67.5,-153</points>
<connection>
<GID>133</GID>
<name>IN_1</name></connection>
<intersection>65.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>77</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>73.5,-142,77.5,-142</points>
<connection>
<GID>129</GID>
<name>OUT</name></connection>
<connection>
<GID>130</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>78</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>83.5,-143,90,-143</points>
<connection>
<GID>130</GID>
<name>OUT</name></connection>
<connection>
<GID>131</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>79</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>95.5,-132.5,110,-132.5</points>
<connection>
<GID>62</GID>
<name>N_in0</name></connection>
<connection>
<GID>126</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>80</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>96,-144,107.5,-144</points>
<connection>
<GID>64</GID>
<name>N_in0</name></connection>
<connection>
<GID>131</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>81</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>96,-154,102.5,-154</points>
<connection>
<GID>66</GID>
<name>N_in0</name></connection>
<connection>
<GID>135</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>82</ID>
<shape>
<hsegment>
<ID>18</ID>
<points>84,-153,90,-153</points>
<connection>
<GID>134</GID>
<name>OUT</name></connection>
<connection>
<GID>135</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>83</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49.5,-150,49.5,-144</points>
<intersection>-150 1</intersection>
<intersection>-144 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>49.5,-150,58.5,-150</points>
<connection>
<GID>132</GID>
<name>IN_0</name></connection>
<intersection>49.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>40.5,-144,49.5,-144</points>
<connection>
<GID>48</GID>
<name>OUT_0</name></connection>
<intersection>49.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>84</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>64.5,-151,67.5,-151</points>
<connection>
<GID>132</GID>
<name>OUT</name></connection>
<connection>
<GID>133</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>85</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73.5,-152,78,-152</points>
<connection>
<GID>133</GID>
<name>OUT</name></connection>
<connection>
<GID>134</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>86</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50.5,-140,50.5,-135.5</points>
<intersection>-140 3</intersection>
<intersection>-135.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>40.5,-135.5,50.5,-135.5</points>
<connection>
<GID>36</GID>
<name>OUT_0</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>50.5,-140,58.5,-140</points>
<connection>
<GID>128</GID>
<name>IN_0</name></connection>
<intersection>50.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>91</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>110,-154,110,-141</points>
<intersection>-154 2</intersection>
<intersection>-141 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>104.5,-154,110,-154</points>
<connection>
<GID>66</GID>
<name>N_in1</name></connection>
<intersection>110 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>110,-141,116,-141</points>
<connection>
<GID>139</GID>
<name>IN_2</name></connection>
<intersection>110 0</intersection></hsegment></shape></wire>
<wire>
<ID>92</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>108.5,-143,108.5,-142</points>
<connection>
<GID>64</GID>
<name>N_in3</name></connection>
<intersection>-142 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>108.5,-142,116,-142</points>
<connection>
<GID>139</GID>
<name>IN_1</name></connection>
<intersection>108.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>93</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>111,-143,111,-133.5</points>
<connection>
<GID>62</GID>
<name>N_in2</name></connection>
<intersection>-143 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>111,-143,116,-143</points>
<connection>
<GID>139</GID>
<name>IN_0</name></connection>
<intersection>111 0</intersection></hsegment></shape></wire>
<wire>
<ID>96</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>92,-104.5,92,-103</points>
<intersection>-104.5 2</intersection>
<intersection>-103 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>92,-103,95.5,-103</points>
<connection>
<GID>142</GID>
<name>IN_0</name></connection>
<intersection>92 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>89,-104.5,92,-104.5</points>
<connection>
<GID>118</GID>
<name>N_in1</name></connection>
<intersection>92 0</intersection></hsegment></shape></wire>
<wire>
<ID>97</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>92,-102,92,-97.5</points>
<intersection>-102 1</intersection>
<intersection>-97.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>92,-102,95.5,-102</points>
<connection>
<GID>142</GID>
<name>IN_1</name></connection>
<intersection>92 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>89,-97.5,92,-97.5</points>
<connection>
<GID>116</GID>
<name>N_in1</name></connection>
<intersection>92 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,4.04748e-006,177.8,-91.7</PageViewport></page 1>
<page 2>
<PageViewport>0,4.04748e-006,177.8,-91.7</PageViewport></page 2>
<page 3>
<PageViewport>0,4.04748e-006,177.8,-91.7</PageViewport></page 3>
<page 4>
<PageViewport>0,4.04748e-006,177.8,-91.7</PageViewport></page 4>
<page 5>
<PageViewport>0,4.04748e-006,177.8,-91.7</PageViewport></page 5>
<page 6>
<PageViewport>0,4.04748e-006,177.8,-91.7</PageViewport></page 6>
<page 7>
<PageViewport>0,4.04748e-006,177.8,-91.7</PageViewport></page 7>
<page 8>
<PageViewport>0,4.04748e-006,177.8,-91.7</PageViewport></page 8>
<page 9>
<PageViewport>0,4.04748e-006,177.8,-91.7</PageViewport></page 9></circuit>