<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>16.0588,-262.364,392.452,-456.488</PageViewport>
<gate>
<ID>1</ID>
<type>AA_LABEL</type>
<position>253.5,-288.5</position>
<gparam>LABEL_TEXT S0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2</ID>
<type>AA_AND2</type>
<position>159,-226</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>3 </input>
<output>
<ID>OUT</ID>4 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3</ID>
<type>AA_LABEL</type>
<position>254.5,-283</position>
<gparam>LABEL_TEXT S1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>4</ID>
<type>AA_AND2</type>
<position>159,-236.5</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>5 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_TOGGLE</type>
<position>123,-225</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>8</ID>
<type>GA_LED</type>
<position>172,-226</position>
<input>
<ID>N_in0</ID>4 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>10</ID>
<type>AA_INVERTER</type>
<position>136,-243.5</position>
<input>
<ID>IN_0</ID>2 </input>
<output>
<ID>OUT_0</ID>3 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>11</ID>
<type>AA_TOGGLE</type>
<position>123,-237</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>12</ID>
<type>GA_LED</type>
<position>172.5,-236.5</position>
<input>
<ID>N_in0</ID>5 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>14</ID>
<type>AA_LABEL</type>
<position>122.5,-222</position>
<gparam>LABEL_TEXT I/p</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>15</ID>
<type>AA_LABEL</type>
<position>119,-234</position>
<gparam>LABEL_TEXT s</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>16</ID>
<type>AA_LABEL</type>
<position>174.5,-222</position>
<gparam>LABEL_TEXT D0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>17</ID>
<type>AA_LABEL</type>
<position>176,-233.5</position>
<gparam>LABEL_TEXT D1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>19</ID>
<type>AA_LABEL</type>
<position>151.5,-214</position>
<gparam>LABEL_TEXT 2x1 De-Multiplexer</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>20</ID>
<type>AA_LABEL</type>
<position>152,-257.5</position>
<gparam>LABEL_TEXT 4x1 De-Multiplexer</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>22</ID>
<type>AA_AND3</type>
<position>162,-280.5</position>
<input>
<ID>IN_0</ID>6 </input>
<input>
<ID>IN_1</ID>9 </input>
<input>
<ID>IN_2</ID>10 </input>
<output>
<ID>OUT</ID>11 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>23</ID>
<type>AA_AND3</type>
<position>162,-289.5</position>
<input>
<ID>IN_0</ID>6 </input>
<input>
<ID>IN_1</ID>9 </input>
<input>
<ID>IN_2</ID>8 </input>
<output>
<ID>OUT</ID>12 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>24</ID>
<type>AA_AND3</type>
<position>162,-298</position>
<input>
<ID>IN_0</ID>6 </input>
<input>
<ID>IN_1</ID>7 </input>
<input>
<ID>IN_2</ID>10 </input>
<output>
<ID>OUT</ID>13 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>25</ID>
<type>AA_AND3</type>
<position>162,-306.5</position>
<input>
<ID>IN_0</ID>6 </input>
<input>
<ID>IN_1</ID>7 </input>
<input>
<ID>IN_2</ID>8 </input>
<output>
<ID>OUT</ID>14 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>27</ID>
<type>AA_TOGGLE</type>
<position>138.5,-266.5</position>
<output>
<ID>OUT_0</ID>8 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>28</ID>
<type>AA_TOGGLE</type>
<position>123.5,-266.5</position>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>29</ID>
<type>AA_TOGGLE</type>
<position>116,-266.5</position>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>31</ID>
<type>AA_LABEL</type>
<position>115,-262.5</position>
<gparam>LABEL_TEXT I/p</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>32</ID>
<type>AA_LABEL</type>
<position>123.5,-262.5</position>
<gparam>LABEL_TEXT S0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>33</ID>
<type>AA_LABEL</type>
<position>138.5,-262.5</position>
<gparam>LABEL_TEXT S1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>35</ID>
<type>AA_INVERTER</type>
<position>144.5,-272</position>
<input>
<ID>IN_0</ID>8 </input>
<output>
<ID>OUT_0</ID>10 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>36</ID>
<type>AA_INVERTER</type>
<position>130,-273.5</position>
<input>
<ID>IN_0</ID>7 </input>
<output>
<ID>OUT_0</ID>9 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>37</ID>
<type>AA_LABEL</type>
<position>166,-274.5</position>
<gparam>LABEL_TEXT D0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>38</ID>
<type>AA_LABEL</type>
<position>166,-284.5</position>
<gparam>LABEL_TEXT D1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>39</ID>
<type>AA_LABEL</type>
<position>167,-293.5</position>
<gparam>LABEL_TEXT D2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>40</ID>
<type>AA_LABEL</type>
<position>167,-302</position>
<gparam>LABEL_TEXT D3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>41</ID>
<type>GA_LED</type>
<position>175.5,-280.5</position>
<input>
<ID>N_in0</ID>11 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>42</ID>
<type>GA_LED</type>
<position>176,-289.5</position>
<input>
<ID>N_in0</ID>12 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>43</ID>
<type>GA_LED</type>
<position>176,-298</position>
<input>
<ID>N_in0</ID>13 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>44</ID>
<type>GA_LED</type>
<position>176.5,-306.5</position>
<input>
<ID>N_in0</ID>14 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>45</ID>
<type>AA_LABEL</type>
<position>138.5,-343.5</position>
<gparam>LABEL_TEXT 8x1 De-Multiplexer</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>47</ID>
<type>AA_TOGGLE</type>
<position>79.5,-366.5</position>
<output>
<ID>OUT_0</ID>15 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>48</ID>
<type>AA_TOGGLE</type>
<position>78.5,-379</position>
<output>
<ID>OUT_0</ID>30 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>49</ID>
<type>AA_TOGGLE</type>
<position>78.5,-396</position>
<output>
<ID>OUT_0</ID>17 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>50</ID>
<type>AA_TOGGLE</type>
<position>79,-413</position>
<output>
<ID>OUT_0</ID>18 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>52</ID>
<type>AA_AND4</type>
<position>130,-359.5</position>
<input>
<ID>IN_0</ID>15 </input>
<input>
<ID>IN_1</ID>19 </input>
<input>
<ID>IN_2</ID>20 </input>
<input>
<ID>IN_3</ID>21 </input>
<output>
<ID>OUT</ID>22 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>54</ID>
<type>AA_AND4</type>
<position>130,-374</position>
<input>
<ID>IN_0</ID>15 </input>
<input>
<ID>IN_1</ID>19 </input>
<input>
<ID>IN_2</ID>20 </input>
<input>
<ID>IN_3</ID>18 </input>
<output>
<ID>OUT</ID>23 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>55</ID>
<type>AA_AND4</type>
<position>130,-388</position>
<input>
<ID>IN_0</ID>15 </input>
<input>
<ID>IN_1</ID>19 </input>
<input>
<ID>IN_2</ID>17 </input>
<input>
<ID>IN_3</ID>21 </input>
<output>
<ID>OUT</ID>24 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>56</ID>
<type>AA_AND4</type>
<position>130,-402</position>
<input>
<ID>IN_0</ID>15 </input>
<input>
<ID>IN_1</ID>19 </input>
<input>
<ID>IN_2</ID>17 </input>
<input>
<ID>IN_3</ID>18 </input>
<output>
<ID>OUT</ID>25 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>57</ID>
<type>AA_AND4</type>
<position>130.5,-416</position>
<input>
<ID>IN_0</ID>15 </input>
<input>
<ID>IN_1</ID>30 </input>
<input>
<ID>IN_2</ID>20 </input>
<input>
<ID>IN_3</ID>21 </input>
<output>
<ID>OUT</ID>26 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>58</ID>
<type>AA_AND4</type>
<position>130.5,-428.5</position>
<input>
<ID>IN_0</ID>15 </input>
<input>
<ID>IN_1</ID>30 </input>
<input>
<ID>IN_2</ID>20 </input>
<input>
<ID>IN_3</ID>18 </input>
<output>
<ID>OUT</ID>27 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>59</ID>
<type>AA_AND4</type>
<position>130.5,-440</position>
<input>
<ID>IN_0</ID>15 </input>
<input>
<ID>IN_1</ID>30 </input>
<input>
<ID>IN_2</ID>17 </input>
<input>
<ID>IN_3</ID>21 </input>
<output>
<ID>OUT</ID>28 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>60</ID>
<type>AA_AND4</type>
<position>130,-452.5</position>
<input>
<ID>IN_0</ID>15 </input>
<input>
<ID>IN_1</ID>30 </input>
<input>
<ID>IN_2</ID>17 </input>
<input>
<ID>IN_3</ID>18 </input>
<output>
<ID>OUT</ID>29 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>62</ID>
<type>AA_LABEL</type>
<position>76,-364.5</position>
<gparam>LABEL_TEXT I/P</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>64</ID>
<type>AA_LABEL</type>
<position>74,-376</position>
<gparam>LABEL_TEXT S0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>65</ID>
<type>AA_LABEL</type>
<position>75,-395</position>
<gparam>LABEL_TEXT S1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>66</ID>
<type>AA_LABEL</type>
<position>74.5,-413</position>
<gparam>LABEL_TEXT S2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>68</ID>
<type>AA_INVERTER</type>
<position>88,-387</position>
<input>
<ID>IN_0</ID>30 </input>
<output>
<ID>OUT_0</ID>19 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>70</ID>
<type>AA_INVERTER</type>
<position>87,-403</position>
<input>
<ID>IN_0</ID>17 </input>
<output>
<ID>OUT_0</ID>20 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>72</ID>
<type>AA_INVERTER</type>
<position>88,-420</position>
<input>
<ID>IN_0</ID>18 </input>
<output>
<ID>OUT_0</ID>21 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>74</ID>
<type>AA_LABEL</type>
<position>135,-352</position>
<gparam>LABEL_TEXT D0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>75</ID>
<type>AA_LABEL</type>
<position>136.5,-369.5</position>
<gparam>LABEL_TEXT D1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>76</ID>
<type>AA_LABEL</type>
<position>136.5,-384</position>
<gparam>LABEL_TEXT D2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>77</ID>
<type>AA_LABEL</type>
<position>137,-397.5</position>
<gparam>LABEL_TEXT D3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>78</ID>
<type>AA_LABEL</type>
<position>136,-411.5</position>
<gparam>LABEL_TEXT D4</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>79</ID>
<type>AA_LABEL</type>
<position>137,-424.5</position>
<gparam>LABEL_TEXT D5</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>80</ID>
<type>AA_LABEL</type>
<position>137,-435.5</position>
<gparam>LABEL_TEXT D6</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>81</ID>
<type>AA_LABEL</type>
<position>137.5,-448</position>
<gparam>LABEL_TEXT D7</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>83</ID>
<type>GA_LED</type>
<position>157.5,-359.5</position>
<input>
<ID>N_in0</ID>22 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>84</ID>
<type>GA_LED</type>
<position>157,-374</position>
<input>
<ID>N_in0</ID>23 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>85</ID>
<type>GA_LED</type>
<position>158,-388</position>
<input>
<ID>N_in0</ID>24 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>86</ID>
<type>GA_LED</type>
<position>158.5,-402</position>
<input>
<ID>N_in0</ID>25 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>87</ID>
<type>GA_LED</type>
<position>157.5,-416</position>
<input>
<ID>N_in0</ID>26 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>88</ID>
<type>GA_LED</type>
<position>158.5,-428.5</position>
<input>
<ID>N_in0</ID>27 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>89</ID>
<type>GA_LED</type>
<position>157.5,-440</position>
<input>
<ID>N_in0</ID>28 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>90</ID>
<type>GA_LED</type>
<position>156.5,-452.5</position>
<input>
<ID>N_in0</ID>29 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>92</ID>
<type>AA_TOGGLE</type>
<position>263,-370</position>
<output>
<ID>OUT_0</ID>31 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>96</ID>
<type>AA_AND4</type>
<position>313.5,-363</position>
<input>
<ID>IN_0</ID>31 </input>
<input>
<ID>IN_1</ID>34 </input>
<input>
<ID>IN_2</ID>35 </input>
<input>
<ID>IN_3</ID>36 </input>
<output>
<ID>OUT</ID>37 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>97</ID>
<type>AA_AND4</type>
<position>313.5,-377.5</position>
<input>
<ID>IN_0</ID>31 </input>
<input>
<ID>IN_1</ID>34 </input>
<input>
<ID>IN_2</ID>35 </input>
<input>
<ID>IN_3</ID>33 </input>
<output>
<ID>OUT</ID>38 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>98</ID>
<type>AA_AND4</type>
<position>313.5,-391.5</position>
<input>
<ID>IN_0</ID>31 </input>
<input>
<ID>IN_1</ID>34 </input>
<input>
<ID>IN_2</ID>32 </input>
<input>
<ID>IN_3</ID>36 </input>
<output>
<ID>OUT</ID>39 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>99</ID>
<type>AA_AND4</type>
<position>313.5,-405.5</position>
<input>
<ID>IN_0</ID>31 </input>
<input>
<ID>IN_1</ID>34 </input>
<input>
<ID>IN_2</ID>32 </input>
<input>
<ID>IN_3</ID>33 </input>
<output>
<ID>OUT</ID>40 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>100</ID>
<type>AA_AND4</type>
<position>314,-419.5</position>
<input>
<ID>IN_0</ID>31 </input>
<input>
<ID>IN_1</ID>45 </input>
<input>
<ID>IN_2</ID>35 </input>
<input>
<ID>IN_3</ID>36 </input>
<output>
<ID>OUT</ID>41 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>101</ID>
<type>AA_AND4</type>
<position>314,-432</position>
<input>
<ID>IN_0</ID>31 </input>
<input>
<ID>IN_1</ID>45 </input>
<input>
<ID>IN_2</ID>35 </input>
<input>
<ID>IN_3</ID>33 </input>
<output>
<ID>OUT</ID>42 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>102</ID>
<type>AA_AND4</type>
<position>314,-443.5</position>
<input>
<ID>IN_0</ID>31 </input>
<input>
<ID>IN_1</ID>45 </input>
<input>
<ID>IN_2</ID>32 </input>
<input>
<ID>IN_3</ID>36 </input>
<output>
<ID>OUT</ID>43 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>103</ID>
<type>AA_AND4</type>
<position>313.5,-456</position>
<input>
<ID>IN_0</ID>31 </input>
<input>
<ID>IN_1</ID>45 </input>
<input>
<ID>IN_2</ID>32 </input>
<input>
<ID>IN_3</ID>33 </input>
<output>
<ID>OUT</ID>44 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>104</ID>
<type>AA_LABEL</type>
<position>259.5,-368</position>
<gparam>LABEL_TEXT I/P</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>105</ID>
<type>AA_LABEL</type>
<position>257.5,-414.5</position>
<gparam>LABEL_TEXT S0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>106</ID>
<type>AA_LABEL</type>
<position>257.5,-397</position>
<gparam>LABEL_TEXT S1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>107</ID>
<type>AA_LABEL</type>
<position>256,-380.5</position>
<gparam>LABEL_TEXT S2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>108</ID>
<type>AA_INVERTER</type>
<position>271.5,-390.5</position>
<input>
<ID>IN_0</ID>45 </input>
<output>
<ID>OUT_0</ID>34 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>109</ID>
<type>AA_INVERTER</type>
<position>270.5,-406.5</position>
<input>
<ID>IN_0</ID>32 </input>
<output>
<ID>OUT_0</ID>35 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>110</ID>
<type>AA_INVERTER</type>
<position>271.5,-423.5</position>
<input>
<ID>IN_0</ID>33 </input>
<output>
<ID>OUT_0</ID>36 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>111</ID>
<type>AA_LABEL</type>
<position>318.5,-355.5</position>
<gparam>LABEL_TEXT D0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>112</ID>
<type>AA_LABEL</type>
<position>320,-373</position>
<gparam>LABEL_TEXT D1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>113</ID>
<type>AA_LABEL</type>
<position>320,-387.5</position>
<gparam>LABEL_TEXT D2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>114</ID>
<type>AA_LABEL</type>
<position>320.5,-401</position>
<gparam>LABEL_TEXT D3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>115</ID>
<type>AA_LABEL</type>
<position>319.5,-415</position>
<gparam>LABEL_TEXT D4</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>116</ID>
<type>AA_LABEL</type>
<position>320.5,-428</position>
<gparam>LABEL_TEXT D5</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>117</ID>
<type>AA_LABEL</type>
<position>320.5,-439</position>
<gparam>LABEL_TEXT D6</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>118</ID>
<type>AA_LABEL</type>
<position>321,-451.5</position>
<gparam>LABEL_TEXT D7</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>119</ID>
<type>GA_LED</type>
<position>341,-363</position>
<input>
<ID>N_in0</ID>37 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>120</ID>
<type>GA_LED</type>
<position>340.5,-377.5</position>
<input>
<ID>N_in0</ID>38 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>121</ID>
<type>GA_LED</type>
<position>341.5,-391.5</position>
<input>
<ID>N_in0</ID>39 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>122</ID>
<type>GA_LED</type>
<position>342,-405.5</position>
<input>
<ID>N_in0</ID>40 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>123</ID>
<type>GA_LED</type>
<position>341,-419.5</position>
<input>
<ID>N_in0</ID>41 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>124</ID>
<type>GA_LED</type>
<position>342,-432</position>
<input>
<ID>N_in0</ID>42 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>125</ID>
<type>GA_LED</type>
<position>341,-443.5</position>
<input>
<ID>N_in0</ID>43 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>126</ID>
<type>GA_LED</type>
<position>340,-456</position>
<input>
<ID>N_in0</ID>44 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>128</ID>
<type>DD_KEYPAD_HEX</type>
<position>220.5,-403.5</position>
<output>
<ID>OUT_0</ID>33 </output>
<output>
<ID>OUT_1</ID>32 </output>
<output>
<ID>OUT_2</ID>45 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>129</ID>
<type>AA_LABEL</type>
<position>298,-260.5</position>
<gparam>LABEL_TEXT 4x1 De-Multiplexer</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>130</ID>
<type>AA_AND3</type>
<position>308,-283.5</position>
<input>
<ID>IN_0</ID>46 </input>
<input>
<ID>IN_1</ID>49 </input>
<input>
<ID>IN_2</ID>50 </input>
<output>
<ID>OUT</ID>51 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>131</ID>
<type>AA_AND3</type>
<position>308,-292.5</position>
<input>
<ID>IN_0</ID>46 </input>
<input>
<ID>IN_1</ID>49 </input>
<input>
<ID>IN_2</ID>48 </input>
<output>
<ID>OUT</ID>52 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>132</ID>
<type>AA_AND3</type>
<position>308,-301</position>
<input>
<ID>IN_0</ID>46 </input>
<input>
<ID>IN_1</ID>47 </input>
<input>
<ID>IN_2</ID>50 </input>
<output>
<ID>OUT</ID>53 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>133</ID>
<type>AA_AND3</type>
<position>308,-309.5</position>
<input>
<ID>IN_0</ID>46 </input>
<input>
<ID>IN_1</ID>47 </input>
<input>
<ID>IN_2</ID>48 </input>
<output>
<ID>OUT</ID>54 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>136</ID>
<type>AA_TOGGLE</type>
<position>262,-269.5</position>
<output>
<ID>OUT_0</ID>46 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>137</ID>
<type>AA_LABEL</type>
<position>261,-265.5</position>
<gparam>LABEL_TEXT I/p</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>140</ID>
<type>AA_INVERTER</type>
<position>290.5,-275</position>
<input>
<ID>IN_0</ID>48 </input>
<output>
<ID>OUT_0</ID>50 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>141</ID>
<type>AA_INVERTER</type>
<position>276,-276.5</position>
<input>
<ID>IN_0</ID>47 </input>
<output>
<ID>OUT_0</ID>49 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>142</ID>
<type>AA_LABEL</type>
<position>312,-277.5</position>
<gparam>LABEL_TEXT D0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>143</ID>
<type>AA_LABEL</type>
<position>312,-287.5</position>
<gparam>LABEL_TEXT D1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>144</ID>
<type>AA_LABEL</type>
<position>313,-296.5</position>
<gparam>LABEL_TEXT D2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>145</ID>
<type>AA_LABEL</type>
<position>313,-305</position>
<gparam>LABEL_TEXT D3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>146</ID>
<type>GA_LED</type>
<position>321.5,-283.5</position>
<input>
<ID>N_in0</ID>51 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>147</ID>
<type>GA_LED</type>
<position>322,-292.5</position>
<input>
<ID>N_in0</ID>52 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>148</ID>
<type>GA_LED</type>
<position>322,-301</position>
<input>
<ID>N_in0</ID>53 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>149</ID>
<type>GA_LED</type>
<position>322.5,-309.5</position>
<input>
<ID>N_in0</ID>54 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>150</ID>
<type>AA_LABEL</type>
<position>298,-344.5</position>
<gparam>LABEL_TEXT 8x1 De-Multiplexer</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>151</ID>
<type>DD_KEYPAD_HEX</type>
<position>244,-284</position>
<output>
<ID>OUT_0</ID>48 </output>
<output>
<ID>OUT_1</ID>47 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<wire>
<ID>1</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>125,-225,156,-225</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<intersection>149.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>149.5,-235.5,149.5,-225</points>
<intersection>-235.5 4</intersection>
<intersection>-225 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>149.5,-235.5,156,-235.5</points>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<intersection>149.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>140.5,-237.5,140.5,-237</points>
<intersection>-237.5 1</intersection>
<intersection>-237 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>140.5,-237.5,156,-237.5</points>
<connection>
<GID>4</GID>
<name>IN_1</name></connection>
<intersection>140.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>125,-237,140.5,-237</points>
<connection>
<GID>11</GID>
<name>OUT_0</name></connection>
<intersection>133 3</intersection>
<intersection>140.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>133,-243.5,133,-237</points>
<connection>
<GID>10</GID>
<name>IN_0</name></connection>
<intersection>-237 2</intersection></vsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>147.5,-243.5,147.5,-227</points>
<intersection>-243.5 2</intersection>
<intersection>-227 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>147.5,-227,156,-227</points>
<connection>
<GID>2</GID>
<name>IN_1</name></connection>
<intersection>147.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>139,-243.5,147.5,-243.5</points>
<connection>
<GID>10</GID>
<name>OUT_0</name></connection>
<intersection>147.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>162,-226,171,-226</points>
<connection>
<GID>2</GID>
<name>OUT</name></connection>
<connection>
<GID>8</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>162,-236.5,171.5,-236.5</points>
<connection>
<GID>4</GID>
<name>OUT</name></connection>
<connection>
<GID>12</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>116,-278.5,116,-268.5</points>
<connection>
<GID>29</GID>
<name>OUT_0</name></connection>
<intersection>-278.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>116,-278.5,159,-278.5</points>
<connection>
<GID>22</GID>
<name>IN_0</name></connection>
<intersection>116 0</intersection>
<intersection>141 2</intersection>
<intersection>150 4</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>141,-304.5,141,-278.5</points>
<intersection>-304.5 3</intersection>
<intersection>-278.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>141,-304.5,159,-304.5</points>
<connection>
<GID>25</GID>
<name>IN_0</name></connection>
<intersection>141 2</intersection>
<intersection>150 6</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>150,-287.5,150,-278.5</points>
<intersection>-287.5 5</intersection>
<intersection>-278.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>150,-287.5,159,-287.5</points>
<connection>
<GID>23</GID>
<name>IN_0</name></connection>
<intersection>150 4</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>150,-304.5,150,-296</points>
<intersection>-304.5 3</intersection>
<intersection>-296 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>150,-296,159,-296</points>
<connection>
<GID>24</GID>
<name>IN_0</name></connection>
<intersection>150 6</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>123.5,-306.5,123.5,-268.5</points>
<connection>
<GID>28</GID>
<name>OUT_0</name></connection>
<intersection>-306.5 1</intersection>
<intersection>-270.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>123.5,-306.5,159,-306.5</points>
<connection>
<GID>25</GID>
<name>IN_1</name></connection>
<intersection>123.5 0</intersection>
<intersection>152.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>123.5,-270.5,130,-270.5</points>
<connection>
<GID>36</GID>
<name>IN_0</name></connection>
<intersection>123.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>152.5,-306.5,152.5,-298</points>
<intersection>-306.5 1</intersection>
<intersection>-298 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>152.5,-298,159,-298</points>
<connection>
<GID>24</GID>
<name>IN_1</name></connection>
<intersection>152.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>138.5,-308.5,138.5,-268.5</points>
<connection>
<GID>27</GID>
<name>OUT_0</name></connection>
<intersection>-308.5 1</intersection>
<intersection>-269 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>138.5,-308.5,159,-308.5</points>
<connection>
<GID>25</GID>
<name>IN_2</name></connection>
<intersection>138.5 0</intersection>
<intersection>147 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>138.5,-269,144.5,-269</points>
<connection>
<GID>35</GID>
<name>IN_0</name></connection>
<intersection>138.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>147,-308.5,147,-291.5</points>
<intersection>-308.5 1</intersection>
<intersection>-291.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>147,-291.5,159,-291.5</points>
<connection>
<GID>23</GID>
<name>IN_2</name></connection>
<intersection>147 3</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>130,-280.5,130,-276.5</points>
<connection>
<GID>36</GID>
<name>OUT_0</name></connection>
<intersection>-280.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>130,-280.5,159,-280.5</points>
<connection>
<GID>22</GID>
<name>IN_1</name></connection>
<intersection>130 0</intersection>
<intersection>156 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>156,-289.5,156,-280.5</points>
<intersection>-289.5 3</intersection>
<intersection>-280.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>156,-289.5,159,-289.5</points>
<connection>
<GID>23</GID>
<name>IN_1</name></connection>
<intersection>156 2</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>144.5,-282.5,144.5,-275</points>
<connection>
<GID>35</GID>
<name>OUT_0</name></connection>
<intersection>-282.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>144.5,-282.5,159,-282.5</points>
<connection>
<GID>22</GID>
<name>IN_2</name></connection>
<intersection>144.5 0</intersection>
<intersection>157 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>157,-300,157,-282.5</points>
<intersection>-300 3</intersection>
<intersection>-282.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>157,-300,159,-300</points>
<connection>
<GID>24</GID>
<name>IN_2</name></connection>
<intersection>157 2</intersection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>165,-280.5,174.5,-280.5</points>
<connection>
<GID>22</GID>
<name>OUT</name></connection>
<connection>
<GID>41</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>165,-289.5,175,-289.5</points>
<connection>
<GID>23</GID>
<name>OUT</name></connection>
<connection>
<GID>42</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>165,-298,175,-298</points>
<connection>
<GID>24</GID>
<name>OUT</name></connection>
<connection>
<GID>43</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>165,-306.5,175.5,-306.5</points>
<connection>
<GID>25</GID>
<name>OUT</name></connection>
<connection>
<GID>44</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>96.5,-449.5,96.5,-356.5</points>
<intersection>-449.5 3</intersection>
<intersection>-366.5 2</intersection>
<intersection>-356.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>96.5,-356.5,127,-356.5</points>
<connection>
<GID>52</GID>
<name>IN_0</name></connection>
<intersection>96.5 0</intersection>
<intersection>122 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>81.5,-366.5,96.5,-366.5</points>
<connection>
<GID>47</GID>
<name>OUT_0</name></connection>
<intersection>96.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>96.5,-449.5,127,-449.5</points>
<connection>
<GID>60</GID>
<name>IN_0</name></connection>
<intersection>96.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>122,-437,122,-356.5</points>
<intersection>-437 16</intersection>
<intersection>-425.5 14</intersection>
<intersection>-413 12</intersection>
<intersection>-399 10</intersection>
<intersection>-385 8</intersection>
<intersection>-371 5</intersection>
<intersection>-356.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>122,-371,127,-371</points>
<connection>
<GID>54</GID>
<name>IN_0</name></connection>
<intersection>122 4</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>122,-385,127,-385</points>
<connection>
<GID>55</GID>
<name>IN_0</name></connection>
<intersection>122 4</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>122,-399,127,-399</points>
<connection>
<GID>56</GID>
<name>IN_0</name></connection>
<intersection>122 4</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>122,-413,127.5,-413</points>
<connection>
<GID>57</GID>
<name>IN_0</name></connection>
<intersection>122 4</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>122,-425.5,127.5,-425.5</points>
<connection>
<GID>58</GID>
<name>IN_0</name></connection>
<intersection>122 4</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>122,-437,127.5,-437</points>
<connection>
<GID>59</GID>
<name>IN_0</name></connection>
<intersection>122 4</intersection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>104,-453.5,104,-396</points>
<intersection>-453.5 1</intersection>
<intersection>-403.5 4</intersection>
<intersection>-396 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>104,-453.5,127,-453.5</points>
<connection>
<GID>60</GID>
<name>IN_2</name></connection>
<intersection>104 0</intersection>
<intersection>126 6</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>80.5,-396,104,-396</points>
<connection>
<GID>49</GID>
<name>OUT_0</name></connection>
<intersection>84 3</intersection>
<intersection>104 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>84,-403,84,-396</points>
<connection>
<GID>70</GID>
<name>IN_0</name></connection>
<intersection>-396 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>104,-403.5,125.5,-403.5</points>
<intersection>104 0</intersection>
<intersection>125.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>125.5,-403.5,125.5,-389</points>
<intersection>-403.5 4</intersection>
<intersection>-403 10</intersection>
<intersection>-389 9</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>126,-453.5,126,-441</points>
<intersection>-453.5 1</intersection>
<intersection>-441 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>126,-441,127.5,-441</points>
<connection>
<GID>59</GID>
<name>IN_2</name></connection>
<intersection>126 6</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>125.5,-389,127,-389</points>
<connection>
<GID>55</GID>
<name>IN_2</name></connection>
<intersection>125.5 5</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>125.5,-403,127,-403</points>
<connection>
<GID>56</GID>
<name>IN_2</name></connection>
<intersection>125.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>101,-455.5,101,-377</points>
<intersection>-455.5 1</intersection>
<intersection>-413 2</intersection>
<intersection>-405 5</intersection>
<intersection>-377 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>101,-455.5,127,-455.5</points>
<connection>
<GID>60</GID>
<name>IN_3</name></connection>
<intersection>101 0</intersection>
<intersection>125 6</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>81,-413,101,-413</points>
<connection>
<GID>50</GID>
<name>OUT_0</name></connection>
<intersection>85 3</intersection>
<intersection>101 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>85,-420,85,-413</points>
<connection>
<GID>72</GID>
<name>IN_0</name></connection>
<intersection>-413 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>101,-377,127,-377</points>
<connection>
<GID>54</GID>
<name>IN_3</name></connection>
<intersection>101 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>101,-405,127,-405</points>
<connection>
<GID>56</GID>
<name>IN_3</name></connection>
<intersection>101 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>125,-455.5,125,-431.5</points>
<intersection>-455.5 1</intersection>
<intersection>-431.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>125,-431.5,127.5,-431.5</points>
<connection>
<GID>58</GID>
<name>IN_3</name></connection>
<intersection>125 6</intersection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>108.5,-387,108.5,-358.5</points>
<intersection>-387 2</intersection>
<intersection>-358.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>108.5,-358.5,127,-358.5</points>
<connection>
<GID>52</GID>
<name>IN_1</name></connection>
<intersection>108.5 0</intersection>
<intersection>124 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>91,-387,108.5,-387</points>
<connection>
<GID>68</GID>
<name>OUT_0</name></connection>
<intersection>108.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>124,-401,124,-358.5</points>
<intersection>-401 9</intersection>
<intersection>-387 7</intersection>
<intersection>-373 5</intersection>
<intersection>-358.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>124,-373,127,-373</points>
<connection>
<GID>54</GID>
<name>IN_1</name></connection>
<intersection>124 4</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>124,-387,127,-387</points>
<connection>
<GID>55</GID>
<name>IN_1</name></connection>
<intersection>124 4</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>124,-401,127,-401</points>
<connection>
<GID>56</GID>
<name>IN_1</name></connection>
<intersection>124 4</intersection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>106.5,-417,106.5,-360.5</points>
<intersection>-417 5</intersection>
<intersection>-403 2</intersection>
<intersection>-360.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>106.5,-360.5,127,-360.5</points>
<connection>
<GID>52</GID>
<name>IN_2</name></connection>
<intersection>106.5 0</intersection>
<intersection>125.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>90,-403,106.5,-403</points>
<connection>
<GID>70</GID>
<name>OUT_0</name></connection>
<intersection>106.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>125.5,-375,125.5,-360.5</points>
<intersection>-375 4</intersection>
<intersection>-360.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>125.5,-375,127,-375</points>
<connection>
<GID>54</GID>
<name>IN_2</name></connection>
<intersection>125.5 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>106.5,-417,127.5,-417</points>
<connection>
<GID>57</GID>
<name>IN_2</name></connection>
<intersection>106.5 0</intersection>
<intersection>125.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>125.5,-429.5,125.5,-417</points>
<intersection>-429.5 7</intersection>
<intersection>-417 5</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>125.5,-429.5,127.5,-429.5</points>
<connection>
<GID>58</GID>
<name>IN_2</name></connection>
<intersection>125.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>110.5,-420,110.5,-362.5</points>
<intersection>-420 2</intersection>
<intersection>-419 4</intersection>
<intersection>-391 3</intersection>
<intersection>-362.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>110.5,-362.5,127,-362.5</points>
<connection>
<GID>52</GID>
<name>IN_3</name></connection>
<intersection>110.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>91,-420,110.5,-420</points>
<connection>
<GID>72</GID>
<name>OUT_0</name></connection>
<intersection>110.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>110.5,-391,127,-391</points>
<connection>
<GID>55</GID>
<name>IN_3</name></connection>
<intersection>110.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>110.5,-419,127.5,-419</points>
<connection>
<GID>57</GID>
<name>IN_3</name></connection>
<intersection>110.5 0</intersection>
<intersection>127 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>127,-443,127,-419</points>
<intersection>-443 6</intersection>
<intersection>-419 4</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>127,-443,127.5,-443</points>
<connection>
<GID>59</GID>
<name>IN_3</name></connection>
<intersection>127 5</intersection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>133,-359.5,156.5,-359.5</points>
<connection>
<GID>52</GID>
<name>OUT</name></connection>
<connection>
<GID>83</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>133,-374,156,-374</points>
<connection>
<GID>54</GID>
<name>OUT</name></connection>
<connection>
<GID>84</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>133,-388,157,-388</points>
<connection>
<GID>55</GID>
<name>OUT</name></connection>
<connection>
<GID>85</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>133,-402,157.5,-402</points>
<connection>
<GID>56</GID>
<name>OUT</name></connection>
<connection>
<GID>86</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>133.5,-416,156.5,-416</points>
<connection>
<GID>57</GID>
<name>OUT</name></connection>
<connection>
<GID>87</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>133.5,-428.5,157.5,-428.5</points>
<connection>
<GID>58</GID>
<name>OUT</name></connection>
<connection>
<GID>88</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>133.5,-440,156.5,-440</points>
<connection>
<GID>59</GID>
<name>OUT</name></connection>
<connection>
<GID>89</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>133,-452.5,155.5,-452.5</points>
<connection>
<GID>60</GID>
<name>OUT</name></connection>
<connection>
<GID>90</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>99,-451.5,99,-379</points>
<intersection>-451.5 1</intersection>
<intersection>-415 4</intersection>
<intersection>-379 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>99,-451.5,127,-451.5</points>
<connection>
<GID>60</GID>
<name>IN_1</name></connection>
<intersection>99 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>80.5,-379,99,-379</points>
<connection>
<GID>48</GID>
<name>OUT_0</name></connection>
<intersection>85 3</intersection>
<intersection>99 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>85,-387,85,-379</points>
<connection>
<GID>68</GID>
<name>IN_0</name></connection>
<intersection>-379 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>99,-415,127.5,-415</points>
<connection>
<GID>57</GID>
<name>IN_1</name></connection>
<intersection>99 0</intersection>
<intersection>123.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>123.5,-439,123.5,-415</points>
<intersection>-439 6</intersection>
<intersection>-427.5 7</intersection>
<intersection>-415 4</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>123.5,-439,127.5,-439</points>
<connection>
<GID>59</GID>
<name>IN_1</name></connection>
<intersection>123.5 5</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>123.5,-427.5,127.5,-427.5</points>
<connection>
<GID>58</GID>
<name>IN_1</name></connection>
<intersection>123.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>280,-453,280,-360</points>
<intersection>-453 3</intersection>
<intersection>-370 2</intersection>
<intersection>-360 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>280,-360,310.5,-360</points>
<connection>
<GID>96</GID>
<name>IN_0</name></connection>
<intersection>280 0</intersection>
<intersection>305.5 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>265,-370,280,-370</points>
<connection>
<GID>92</GID>
<name>OUT_0</name></connection>
<intersection>280 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>280,-453,310.5,-453</points>
<connection>
<GID>103</GID>
<name>IN_0</name></connection>
<intersection>280 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>305.5,-440.5,305.5,-360</points>
<intersection>-440.5 16</intersection>
<intersection>-429 14</intersection>
<intersection>-416.5 12</intersection>
<intersection>-402.5 10</intersection>
<intersection>-388.5 8</intersection>
<intersection>-374.5 5</intersection>
<intersection>-360 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>305.5,-374.5,310.5,-374.5</points>
<connection>
<GID>97</GID>
<name>IN_0</name></connection>
<intersection>305.5 4</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>305.5,-388.5,310.5,-388.5</points>
<connection>
<GID>98</GID>
<name>IN_0</name></connection>
<intersection>305.5 4</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>305.5,-402.5,310.5,-402.5</points>
<connection>
<GID>99</GID>
<name>IN_0</name></connection>
<intersection>305.5 4</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>305.5,-416.5,311,-416.5</points>
<connection>
<GID>100</GID>
<name>IN_0</name></connection>
<intersection>305.5 4</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>305.5,-429,311,-429</points>
<connection>
<GID>101</GID>
<name>IN_0</name></connection>
<intersection>305.5 4</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>305.5,-440.5,311,-440.5</points>
<connection>
<GID>102</GID>
<name>IN_0</name></connection>
<intersection>305.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>287.5,-457,287.5,-399.5</points>
<intersection>-457 1</intersection>
<intersection>-407 4</intersection>
<intersection>-399.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>287.5,-457,310.5,-457</points>
<connection>
<GID>103</GID>
<name>IN_2</name></connection>
<intersection>287.5 0</intersection>
<intersection>309.5 6</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>237,-399.5,287.5,-399.5</points>
<intersection>237 12</intersection>
<intersection>267.5 3</intersection>
<intersection>287.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>267.5,-406.5,267.5,-399.5</points>
<connection>
<GID>109</GID>
<name>IN_0</name></connection>
<intersection>-399.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>287.5,-407,309,-407</points>
<intersection>287.5 0</intersection>
<intersection>309 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>309,-407,309,-392.5</points>
<intersection>-407 4</intersection>
<intersection>-406.5 10</intersection>
<intersection>-392.5 9</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>309.5,-457,309.5,-444.5</points>
<intersection>-457 1</intersection>
<intersection>-444.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>309.5,-444.5,311,-444.5</points>
<connection>
<GID>102</GID>
<name>IN_2</name></connection>
<intersection>309.5 6</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>309,-392.5,310.5,-392.5</points>
<connection>
<GID>98</GID>
<name>IN_2</name></connection>
<intersection>309 5</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>309,-406.5,310.5,-406.5</points>
<connection>
<GID>99</GID>
<name>IN_2</name></connection>
<intersection>309 5</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>237,-404.5,237,-399.5</points>
<intersection>-404.5 13</intersection>
<intersection>-399.5 2</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>225.5,-404.5,237,-404.5</points>
<connection>
<GID>128</GID>
<name>OUT_1</name></connection>
<intersection>237 12</intersection></hsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>284.5,-459,284.5,-380.5</points>
<intersection>-459 1</intersection>
<intersection>-416.5 2</intersection>
<intersection>-408.5 5</intersection>
<intersection>-380.5 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>284.5,-459,310.5,-459</points>
<connection>
<GID>103</GID>
<name>IN_3</name></connection>
<intersection>284.5 0</intersection>
<intersection>308.5 6</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>225.5,-416.5,284.5,-416.5</points>
<intersection>225.5 9</intersection>
<intersection>268.5 3</intersection>
<intersection>284.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>268.5,-423.5,268.5,-416.5</points>
<connection>
<GID>110</GID>
<name>IN_0</name></connection>
<intersection>-416.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>284.5,-380.5,310.5,-380.5</points>
<connection>
<GID>97</GID>
<name>IN_3</name></connection>
<intersection>284.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>284.5,-408.5,310.5,-408.5</points>
<connection>
<GID>99</GID>
<name>IN_3</name></connection>
<intersection>284.5 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>308.5,-459,308.5,-435</points>
<intersection>-459 1</intersection>
<intersection>-435 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>308.5,-435,311,-435</points>
<connection>
<GID>101</GID>
<name>IN_3</name></connection>
<intersection>308.5 6</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>225.5,-416.5,225.5,-406.5</points>
<connection>
<GID>128</GID>
<name>OUT_0</name></connection>
<intersection>-416.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>292,-390.5,292,-362</points>
<intersection>-390.5 2</intersection>
<intersection>-362 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>292,-362,310.5,-362</points>
<connection>
<GID>96</GID>
<name>IN_1</name></connection>
<intersection>292 0</intersection>
<intersection>307.5 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>274.5,-390.5,310.5,-390.5</points>
<connection>
<GID>98</GID>
<name>IN_1</name></connection>
<connection>
<GID>108</GID>
<name>OUT_0</name></connection>
<intersection>292 0</intersection>
<intersection>307.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>307.5,-404.5,307.5,-362</points>
<intersection>-404.5 9</intersection>
<intersection>-390.5 2</intersection>
<intersection>-376.5 5</intersection>
<intersection>-362 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>307.5,-376.5,310.5,-376.5</points>
<connection>
<GID>97</GID>
<name>IN_1</name></connection>
<intersection>307.5 4</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>307.5,-404.5,310.5,-404.5</points>
<connection>
<GID>99</GID>
<name>IN_1</name></connection>
<intersection>307.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>290,-433,290,-364</points>
<intersection>-433 5</intersection>
<intersection>-406.5 2</intersection>
<intersection>-364 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>290,-364,310.5,-364</points>
<connection>
<GID>96</GID>
<name>IN_2</name></connection>
<intersection>290 0</intersection>
<intersection>309 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>273.5,-406.5,290,-406.5</points>
<connection>
<GID>109</GID>
<name>OUT_0</name></connection>
<intersection>290 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>309,-378.5,309,-364</points>
<intersection>-378.5 4</intersection>
<intersection>-364 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>309,-378.5,310.5,-378.5</points>
<connection>
<GID>97</GID>
<name>IN_2</name></connection>
<intersection>309 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>290,-433,311,-433</points>
<connection>
<GID>101</GID>
<name>IN_2</name></connection>
<intersection>290 0</intersection>
<intersection>311 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>311,-433,311,-420.5</points>
<connection>
<GID>100</GID>
<name>IN_2</name></connection>
<intersection>-433 5</intersection></vsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>294,-423.5,294,-366</points>
<intersection>-423.5 2</intersection>
<intersection>-422.5 4</intersection>
<intersection>-394.5 3</intersection>
<intersection>-366 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>294,-366,310.5,-366</points>
<connection>
<GID>96</GID>
<name>IN_3</name></connection>
<intersection>294 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>274.5,-423.5,294,-423.5</points>
<connection>
<GID>110</GID>
<name>OUT_0</name></connection>
<intersection>294 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>294,-394.5,310.5,-394.5</points>
<connection>
<GID>98</GID>
<name>IN_3</name></connection>
<intersection>294 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>294,-422.5,311,-422.5</points>
<connection>
<GID>100</GID>
<name>IN_3</name></connection>
<intersection>294 0</intersection>
<intersection>310.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>310.5,-446.5,310.5,-422.5</points>
<intersection>-446.5 6</intersection>
<intersection>-422.5 4</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>310.5,-446.5,311,-446.5</points>
<connection>
<GID>102</GID>
<name>IN_3</name></connection>
<intersection>310.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>316.5,-363,340,-363</points>
<connection>
<GID>96</GID>
<name>OUT</name></connection>
<connection>
<GID>119</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>316.5,-377.5,339.5,-377.5</points>
<connection>
<GID>97</GID>
<name>OUT</name></connection>
<connection>
<GID>120</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>316.5,-391.5,340.5,-391.5</points>
<connection>
<GID>98</GID>
<name>OUT</name></connection>
<connection>
<GID>121</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>316.5,-405.5,341,-405.5</points>
<connection>
<GID>99</GID>
<name>OUT</name></connection>
<connection>
<GID>122</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>317,-419.5,340,-419.5</points>
<connection>
<GID>100</GID>
<name>OUT</name></connection>
<connection>
<GID>123</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>317,-432,341,-432</points>
<connection>
<GID>101</GID>
<name>OUT</name></connection>
<connection>
<GID>124</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>317,-443.5,340,-443.5</points>
<connection>
<GID>102</GID>
<name>OUT</name></connection>
<connection>
<GID>125</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>316.5,-456,339,-456</points>
<connection>
<GID>103</GID>
<name>OUT</name></connection>
<connection>
<GID>126</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>282.5,-455,282.5,-382.5</points>
<intersection>-455 1</intersection>
<intersection>-418.5 4</intersection>
<intersection>-382.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>282.5,-455,310.5,-455</points>
<connection>
<GID>103</GID>
<name>IN_1</name></connection>
<intersection>282.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>225.5,-382.5,282.5,-382.5</points>
<intersection>225.5 9</intersection>
<intersection>268.5 3</intersection>
<intersection>282.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>268.5,-390.5,268.5,-382.5</points>
<connection>
<GID>108</GID>
<name>IN_0</name></connection>
<intersection>-382.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>282.5,-418.5,311,-418.5</points>
<connection>
<GID>100</GID>
<name>IN_1</name></connection>
<intersection>282.5 0</intersection>
<intersection>307 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>307,-442.5,307,-418.5</points>
<intersection>-442.5 6</intersection>
<intersection>-431 7</intersection>
<intersection>-418.5 4</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>307,-442.5,311,-442.5</points>
<connection>
<GID>102</GID>
<name>IN_1</name></connection>
<intersection>307 5</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>307,-431,311,-431</points>
<connection>
<GID>101</GID>
<name>IN_1</name></connection>
<intersection>307 5</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>225.5,-402.5,225.5,-382.5</points>
<connection>
<GID>128</GID>
<name>OUT_2</name></connection>
<intersection>-382.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>46</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>262,-281.5,262,-271.5</points>
<connection>
<GID>136</GID>
<name>OUT_0</name></connection>
<intersection>-281.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>262,-281.5,305,-281.5</points>
<connection>
<GID>130</GID>
<name>IN_0</name></connection>
<intersection>262 0</intersection>
<intersection>287 2</intersection>
<intersection>296 4</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>287,-307.5,287,-281.5</points>
<intersection>-307.5 3</intersection>
<intersection>-281.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>287,-307.5,305,-307.5</points>
<connection>
<GID>133</GID>
<name>IN_0</name></connection>
<intersection>287 2</intersection>
<intersection>296 6</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>296,-290.5,296,-281.5</points>
<intersection>-290.5 5</intersection>
<intersection>-281.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>296,-290.5,305,-290.5</points>
<connection>
<GID>131</GID>
<name>IN_0</name></connection>
<intersection>296 4</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>296,-307.5,296,-299</points>
<intersection>-307.5 3</intersection>
<intersection>-299 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>296,-299,305,-299</points>
<connection>
<GID>132</GID>
<name>IN_0</name></connection>
<intersection>296 6</intersection></hsegment></shape></wire>
<wire>
<ID>47</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>269.5,-309.5,269.5,-273.5</points>
<intersection>-309.5 1</intersection>
<intersection>-285 8</intersection>
<intersection>-273.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>269.5,-309.5,305,-309.5</points>
<connection>
<GID>133</GID>
<name>IN_1</name></connection>
<intersection>269.5 0</intersection>
<intersection>298.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>269.5,-273.5,276,-273.5</points>
<connection>
<GID>141</GID>
<name>IN_0</name></connection>
<intersection>269.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>298.5,-309.5,298.5,-301</points>
<intersection>-309.5 1</intersection>
<intersection>-301 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>298.5,-301,305,-301</points>
<connection>
<GID>132</GID>
<name>IN_1</name></connection>
<intersection>298.5 3</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>249,-285,269.5,-285</points>
<connection>
<GID>151</GID>
<name>OUT_1</name></connection>
<intersection>269.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>284.5,-311.5,284.5,-272</points>
<intersection>-311.5 1</intersection>
<intersection>-287 8</intersection>
<intersection>-272 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>284.5,-311.5,305,-311.5</points>
<connection>
<GID>133</GID>
<name>IN_2</name></connection>
<intersection>284.5 0</intersection>
<intersection>293 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>284.5,-272,290.5,-272</points>
<connection>
<GID>140</GID>
<name>IN_0</name></connection>
<intersection>284.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>293,-311.5,293,-294.5</points>
<intersection>-311.5 1</intersection>
<intersection>-294.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>293,-294.5,305,-294.5</points>
<connection>
<GID>131</GID>
<name>IN_2</name></connection>
<intersection>293 3</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>249,-287,284.5,-287</points>
<connection>
<GID>151</GID>
<name>OUT_0</name></connection>
<intersection>284.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>276,-283.5,276,-279.5</points>
<connection>
<GID>141</GID>
<name>OUT_0</name></connection>
<intersection>-283.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>276,-283.5,305,-283.5</points>
<connection>
<GID>130</GID>
<name>IN_1</name></connection>
<intersection>276 0</intersection>
<intersection>302 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>302,-292.5,302,-283.5</points>
<intersection>-292.5 3</intersection>
<intersection>-283.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>302,-292.5,305,-292.5</points>
<connection>
<GID>131</GID>
<name>IN_1</name></connection>
<intersection>302 2</intersection></hsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>290.5,-285.5,290.5,-278</points>
<connection>
<GID>140</GID>
<name>OUT_0</name></connection>
<intersection>-285.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>290.5,-285.5,305,-285.5</points>
<connection>
<GID>130</GID>
<name>IN_2</name></connection>
<intersection>290.5 0</intersection>
<intersection>303 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>303,-303,303,-285.5</points>
<intersection>-303 3</intersection>
<intersection>-285.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>303,-303,305,-303</points>
<connection>
<GID>132</GID>
<name>IN_2</name></connection>
<intersection>303 2</intersection></hsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>311,-283.5,320.5,-283.5</points>
<connection>
<GID>146</GID>
<name>N_in0</name></connection>
<connection>
<GID>130</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>52</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>311,-292.5,321,-292.5</points>
<connection>
<GID>147</GID>
<name>N_in0</name></connection>
<connection>
<GID>131</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>53</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>311,-301,321,-301</points>
<connection>
<GID>148</GID>
<name>N_in0</name></connection>
<connection>
<GID>132</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>54</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>311,-309.5,321.5,-309.5</points>
<connection>
<GID>149</GID>
<name>N_in0</name></connection>
<connection>
<GID>133</GID>
<name>OUT</name></connection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,46.8717,715.223,-322.003</PageViewport></page 1>
<page 2>
<PageViewport>0,46.8717,715.223,-322.003</PageViewport></page 2>
<page 3>
<PageViewport>0,46.8717,715.223,-322.003</PageViewport></page 3>
<page 4>
<PageViewport>0,46.8717,715.223,-322.003</PageViewport></page 4>
<page 5>
<PageViewport>0,46.8717,715.223,-322.003</PageViewport></page 5>
<page 6>
<PageViewport>0,46.8717,715.223,-322.003</PageViewport></page 6>
<page 7>
<PageViewport>0,46.8717,715.223,-322.003</PageViewport></page 7>
<page 8>
<PageViewport>0,46.8717,715.223,-322.003</PageViewport></page 8>
<page 9>
<PageViewport>0,46.8717,715.223,-322.003</PageViewport></page 9></circuit>