<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-98.1295,2.05824,388.158,-248.744</PageViewport>
<gate>
<ID>2</ID>
<type>BA_NAND2</type>
<position>54,-28</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>3 </input>
<output>
<ID>OUT</ID>4 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3</ID>
<type>BA_NAND2</type>
<position>53.5,-42</position>
<input>
<ID>IN_0</ID>3 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>5 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4</ID>
<type>BA_NAND2</type>
<position>75,-29</position>
<input>
<ID>IN_0</ID>4 </input>
<input>
<ID>IN_1</ID>6 </input>
<output>
<ID>OUT</ID>7 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5</ID>
<type>BA_NAND2</type>
<position>75,-39.5</position>
<input>
<ID>IN_0</ID>7 </input>
<input>
<ID>IN_1</ID>5 </input>
<output>
<ID>OUT</ID>6 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7</ID>
<type>AA_INVERTER</type>
<position>38,-34.5</position>
<input>
<ID>IN_0</ID>1 </input>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>9</ID>
<type>AA_TOGGLE</type>
<position>27,-27</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>11</ID>
<type>GA_LED</type>
<position>93,-29</position>
<input>
<ID>N_in0</ID>7 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>13</ID>
<type>GA_LED</type>
<position>92.5,-39.5</position>
<input>
<ID>N_in0</ID>6 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>15</ID>
<type>AA_TOGGLE</type>
<position>42.5,-35</position>
<output>
<ID>OUT_0</ID>3 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>17</ID>
<type>AA_LABEL</type>
<position>25.5,-22.5</position>
<gparam>LABEL_TEXT D</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>18</ID>
<type>AA_LABEL</type>
<position>93,-24</position>
<gparam>LABEL_TEXT Q</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>19</ID>
<type>AA_LABEL</type>
<position>93.5,-36</position>
<gparam>LABEL_TEXT Q`</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>20</ID>
<type>AA_LABEL</type>
<position>42,-31</position>
<gparam>LABEL_TEXT En</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>21</ID>
<type>BA_NAND2</type>
<position>50.5,-71</position>
<input>
<ID>IN_0</ID>8 </input>
<input>
<ID>IN_1</ID>10 </input>
<output>
<ID>OUT</ID>11 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>22</ID>
<type>BA_NAND2</type>
<position>50,-82.5</position>
<input>
<ID>IN_0</ID>10 </input>
<input>
<ID>IN_1</ID>9 </input>
<output>
<ID>OUT</ID>12 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>23</ID>
<type>BA_NAND2</type>
<position>71.5,-72</position>
<input>
<ID>IN_0</ID>11 </input>
<input>
<ID>IN_1</ID>13 </input>
<output>
<ID>OUT</ID>14 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>24</ID>
<type>BA_NAND2</type>
<position>71.5,-80</position>
<input>
<ID>IN_0</ID>14 </input>
<input>
<ID>IN_1</ID>12 </input>
<output>
<ID>OUT</ID>13 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>25</ID>
<type>AA_INVERTER</type>
<position>32.5,-77</position>
<input>
<ID>IN_0</ID>8 </input>
<output>
<ID>OUT_0</ID>9 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>27</ID>
<type>GA_LED</type>
<position>89.5,-72</position>
<input>
<ID>N_in0</ID>14 </input>
<input>
<ID>N_in1</ID>99 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>28</ID>
<type>GA_LED</type>
<position>89,-80</position>
<input>
<ID>N_in0</ID>13 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>31</ID>
<type>AA_LABEL</type>
<position>89.5,-67</position>
<gparam>LABEL_TEXT Q</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>32</ID>
<type>AA_LABEL</type>
<position>90,-76.5</position>
<gparam>LABEL_TEXT Q`</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>35</ID>
<type>BB_CLOCK</type>
<position>38.5,-75</position>
<output>
<ID>CLK</ID>10 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>36</ID>
<type>BA_NAND2</type>
<position>49,-89</position>
<input>
<ID>IN_0</ID>15 </input>
<input>
<ID>IN_1</ID>17 </input>
<output>
<ID>OUT</ID>18 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>37</ID>
<type>BA_NAND2</type>
<position>48.5,-103</position>
<input>
<ID>IN_0</ID>17 </input>
<input>
<ID>IN_1</ID>16 </input>
<output>
<ID>OUT</ID>19 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>38</ID>
<type>BA_NAND2</type>
<position>70,-90</position>
<input>
<ID>IN_0</ID>18 </input>
<input>
<ID>IN_1</ID>20 </input>
<output>
<ID>OUT</ID>21 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>39</ID>
<type>BA_NAND2</type>
<position>70,-100.5</position>
<input>
<ID>IN_0</ID>21 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>20 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>40</ID>
<type>AA_INVERTER</type>
<position>31,-95</position>
<input>
<ID>IN_0</ID>15 </input>
<output>
<ID>OUT_0</ID>16 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>42</ID>
<type>GA_LED</type>
<position>88,-90</position>
<input>
<ID>N_in0</ID>21 </input>
<input>
<ID>N_in1</ID>100 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>43</ID>
<type>GA_LED</type>
<position>87.5,-100.5</position>
<input>
<ID>N_in0</ID>20 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>45</ID>
<type>AA_LABEL</type>
<position>88,-85</position>
<gparam>LABEL_TEXT Q</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>46</ID>
<type>AA_LABEL</type>
<position>88.5,-97</position>
<gparam>LABEL_TEXT Q`</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>47</ID>
<type>BB_CLOCK</type>
<position>37,-95.5</position>
<output>
<ID>CLK</ID>17 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>48</ID>
<type>BA_NAND2</type>
<position>49.5,-111</position>
<input>
<ID>IN_0</ID>22 </input>
<input>
<ID>IN_1</ID>24 </input>
<output>
<ID>OUT</ID>25 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>49</ID>
<type>BA_NAND2</type>
<position>49,-125</position>
<input>
<ID>IN_0</ID>24 </input>
<input>
<ID>IN_1</ID>23 </input>
<output>
<ID>OUT</ID>26 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>50</ID>
<type>BA_NAND2</type>
<position>70.5,-112</position>
<input>
<ID>IN_0</ID>25 </input>
<input>
<ID>IN_1</ID>27 </input>
<output>
<ID>OUT</ID>28 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>51</ID>
<type>BA_NAND2</type>
<position>70.5,-122.5</position>
<input>
<ID>IN_0</ID>28 </input>
<input>
<ID>IN_1</ID>26 </input>
<output>
<ID>OUT</ID>27 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>52</ID>
<type>AA_INVERTER</type>
<position>31.5,-117</position>
<input>
<ID>IN_0</ID>22 </input>
<output>
<ID>OUT_0</ID>23 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>54</ID>
<type>GA_LED</type>
<position>88.5,-112</position>
<input>
<ID>N_in0</ID>28 </input>
<input>
<ID>N_in1</ID>101 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>55</ID>
<type>GA_LED</type>
<position>88,-122.5</position>
<input>
<ID>N_in0</ID>27 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>57</ID>
<type>AA_LABEL</type>
<position>88.5,-107</position>
<gparam>LABEL_TEXT Q</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>58</ID>
<type>AA_LABEL</type>
<position>89,-119</position>
<gparam>LABEL_TEXT Q`</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>59</ID>
<type>BB_CLOCK</type>
<position>37.5,-117.5</position>
<output>
<ID>CLK</ID>24 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>60</ID>
<type>BA_NAND2</type>
<position>50.5,-133.5</position>
<input>
<ID>IN_0</ID>29 </input>
<input>
<ID>IN_1</ID>31 </input>
<output>
<ID>OUT</ID>32 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>61</ID>
<type>BA_NAND2</type>
<position>50,-147.5</position>
<input>
<ID>IN_0</ID>31 </input>
<input>
<ID>IN_1</ID>30 </input>
<output>
<ID>OUT</ID>33 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>62</ID>
<type>BA_NAND2</type>
<position>71.5,-134.5</position>
<input>
<ID>IN_0</ID>32 </input>
<input>
<ID>IN_1</ID>34 </input>
<output>
<ID>OUT</ID>35 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>63</ID>
<type>BA_NAND2</type>
<position>71.5,-145</position>
<input>
<ID>IN_0</ID>35 </input>
<input>
<ID>IN_1</ID>33 </input>
<output>
<ID>OUT</ID>34 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>64</ID>
<type>AA_INVERTER</type>
<position>32.5,-139.5</position>
<input>
<ID>IN_0</ID>29 </input>
<output>
<ID>OUT_0</ID>30 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>66</ID>
<type>GA_LED</type>
<position>89.5,-134.5</position>
<input>
<ID>N_in0</ID>35 </input>
<input>
<ID>N_in1</ID>102 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>67</ID>
<type>GA_LED</type>
<position>89,-145</position>
<input>
<ID>N_in0</ID>34 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>69</ID>
<type>AA_LABEL</type>
<position>89.5,-129.5</position>
<gparam>LABEL_TEXT Q</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>70</ID>
<type>AA_LABEL</type>
<position>90,-141.5</position>
<gparam>LABEL_TEXT Q`</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>71</ID>
<type>BB_CLOCK</type>
<position>38.5,-140</position>
<output>
<ID>CLK</ID>31 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>123</ID>
<type>DD_KEYPAD_HEX</type>
<position>-42.5,-133</position>
<output>
<ID>OUT_0</ID>8 </output>
<output>
<ID>OUT_1</ID>15 </output>
<output>
<ID>OUT_2</ID>22 </output>
<output>
<ID>OUT_3</ID>29 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 10</lparam></gate>
<gate>
<ID>136</ID>
<type>BA_NAND2</type>
<position>50.5,-158.5</position>
<input>
<ID>IN_0</ID>71 </input>
<input>
<ID>IN_1</ID>73 </input>
<output>
<ID>OUT</ID>74 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>137</ID>
<type>BA_NAND2</type>
<position>50,-170</position>
<input>
<ID>IN_0</ID>73 </input>
<input>
<ID>IN_1</ID>72 </input>
<output>
<ID>OUT</ID>75 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>138</ID>
<type>BA_NAND2</type>
<position>71.5,-159.5</position>
<input>
<ID>IN_0</ID>74 </input>
<input>
<ID>IN_1</ID>76 </input>
<output>
<ID>OUT</ID>77 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>139</ID>
<type>BA_NAND2</type>
<position>71.5,-167.5</position>
<input>
<ID>IN_0</ID>77 </input>
<input>
<ID>IN_1</ID>75 </input>
<output>
<ID>OUT</ID>76 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>140</ID>
<type>AA_INVERTER</type>
<position>32.5,-164.5</position>
<input>
<ID>IN_0</ID>71 </input>
<output>
<ID>OUT_0</ID>72 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>141</ID>
<type>GA_LED</type>
<position>89.5,-159.5</position>
<input>
<ID>N_in0</ID>77 </input>
<input>
<ID>N_in1</ID>103 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>142</ID>
<type>GA_LED</type>
<position>89,-167.5</position>
<input>
<ID>N_in0</ID>76 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>143</ID>
<type>AA_LABEL</type>
<position>89.5,-154.5</position>
<gparam>LABEL_TEXT Q</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>144</ID>
<type>AA_LABEL</type>
<position>90,-164</position>
<gparam>LABEL_TEXT Q`</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>145</ID>
<type>BB_CLOCK</type>
<position>38.5,-162.5</position>
<output>
<ID>CLK</ID>73 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>146</ID>
<type>BA_NAND2</type>
<position>49,-176.5</position>
<input>
<ID>IN_0</ID>78 </input>
<input>
<ID>IN_1</ID>80 </input>
<output>
<ID>OUT</ID>81 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>147</ID>
<type>BA_NAND2</type>
<position>48.5,-190.5</position>
<input>
<ID>IN_0</ID>80 </input>
<input>
<ID>IN_1</ID>79 </input>
<output>
<ID>OUT</ID>82 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>148</ID>
<type>BA_NAND2</type>
<position>70,-177.5</position>
<input>
<ID>IN_0</ID>81 </input>
<input>
<ID>IN_1</ID>83 </input>
<output>
<ID>OUT</ID>84 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>149</ID>
<type>BA_NAND2</type>
<position>70,-188</position>
<input>
<ID>IN_0</ID>84 </input>
<input>
<ID>IN_1</ID>82 </input>
<output>
<ID>OUT</ID>83 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>150</ID>
<type>AA_INVERTER</type>
<position>31,-182.5</position>
<input>
<ID>IN_0</ID>78 </input>
<output>
<ID>OUT_0</ID>79 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>151</ID>
<type>GA_LED</type>
<position>88,-177.5</position>
<input>
<ID>N_in0</ID>84 </input>
<input>
<ID>N_in1</ID>104 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>152</ID>
<type>GA_LED</type>
<position>87.5,-188</position>
<input>
<ID>N_in0</ID>83 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>153</ID>
<type>AA_LABEL</type>
<position>88,-172.5</position>
<gparam>LABEL_TEXT Q</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>154</ID>
<type>AA_LABEL</type>
<position>88.5,-184.5</position>
<gparam>LABEL_TEXT Q`</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>155</ID>
<type>BB_CLOCK</type>
<position>37,-183</position>
<output>
<ID>CLK</ID>80 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>156</ID>
<type>BA_NAND2</type>
<position>49.5,-198.5</position>
<input>
<ID>IN_0</ID>85 </input>
<input>
<ID>IN_1</ID>87 </input>
<output>
<ID>OUT</ID>88 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>157</ID>
<type>BA_NAND2</type>
<position>49,-212.5</position>
<input>
<ID>IN_0</ID>87 </input>
<input>
<ID>IN_1</ID>86 </input>
<output>
<ID>OUT</ID>89 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>158</ID>
<type>BA_NAND2</type>
<position>70.5,-199.5</position>
<input>
<ID>IN_0</ID>88 </input>
<input>
<ID>IN_1</ID>90 </input>
<output>
<ID>OUT</ID>91 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>159</ID>
<type>BA_NAND2</type>
<position>70.5,-210</position>
<input>
<ID>IN_0</ID>91 </input>
<input>
<ID>IN_1</ID>89 </input>
<output>
<ID>OUT</ID>90 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>160</ID>
<type>AA_INVERTER</type>
<position>31.5,-204.5</position>
<input>
<ID>IN_0</ID>85 </input>
<output>
<ID>OUT_0</ID>86 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>161</ID>
<type>GA_LED</type>
<position>88.5,-199.5</position>
<input>
<ID>N_in0</ID>91 </input>
<input>
<ID>N_in1</ID>105 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>162</ID>
<type>GA_LED</type>
<position>88,-210</position>
<input>
<ID>N_in0</ID>90 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>163</ID>
<type>AA_LABEL</type>
<position>88.5,-194.5</position>
<gparam>LABEL_TEXT Q</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>164</ID>
<type>AA_LABEL</type>
<position>89,-206.5</position>
<gparam>LABEL_TEXT Q`</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>165</ID>
<type>BB_CLOCK</type>
<position>37.5,-205</position>
<output>
<ID>CLK</ID>87 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>166</ID>
<type>BA_NAND2</type>
<position>50.5,-221</position>
<input>
<ID>IN_0</ID>92 </input>
<input>
<ID>IN_1</ID>94 </input>
<output>
<ID>OUT</ID>95 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>167</ID>
<type>BA_NAND2</type>
<position>50,-235</position>
<input>
<ID>IN_0</ID>94 </input>
<input>
<ID>IN_1</ID>93 </input>
<output>
<ID>OUT</ID>96 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>168</ID>
<type>BA_NAND2</type>
<position>71.5,-222</position>
<input>
<ID>IN_0</ID>95 </input>
<input>
<ID>IN_1</ID>97 </input>
<output>
<ID>OUT</ID>98 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>169</ID>
<type>BA_NAND2</type>
<position>71.5,-232.5</position>
<input>
<ID>IN_0</ID>98 </input>
<input>
<ID>IN_1</ID>96 </input>
<output>
<ID>OUT</ID>97 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>170</ID>
<type>AA_INVERTER</type>
<position>32.5,-227</position>
<input>
<ID>IN_0</ID>92 </input>
<output>
<ID>OUT_0</ID>93 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>171</ID>
<type>GA_LED</type>
<position>89.5,-222</position>
<input>
<ID>N_in0</ID>98 </input>
<input>
<ID>N_in1</ID>106 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>172</ID>
<type>GA_LED</type>
<position>89,-232.5</position>
<input>
<ID>N_in0</ID>97 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>173</ID>
<type>AA_LABEL</type>
<position>89.5,-217</position>
<gparam>LABEL_TEXT Q</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>174</ID>
<type>AA_LABEL</type>
<position>90,-229</position>
<gparam>LABEL_TEXT Q`</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>175</ID>
<type>BB_CLOCK</type>
<position>38.5,-227.5</position>
<output>
<ID>CLK</ID>94 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>176</ID>
<type>DD_KEYPAD_HEX</type>
<position>-43,-152</position>
<output>
<ID>OUT_0</ID>71 </output>
<output>
<ID>OUT_1</ID>78 </output>
<output>
<ID>OUT_2</ID>85 </output>
<output>
<ID>OUT_3</ID>92 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 10</lparam></gate>
<gate>
<ID>178</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>164,-144</position>
<input>
<ID>IN_0</ID>99 </input>
<input>
<ID>IN_1</ID>100 </input>
<input>
<ID>IN_2</ID>101 </input>
<input>
<ID>IN_3</ID>102 </input>
<input>
<ID>IN_4</ID>103 </input>
<input>
<ID>IN_5</ID>104 </input>
<input>
<ID>IN_6</ID>105 </input>
<input>
<ID>IN_7</ID>106 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 170</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<wire>
<ID>1</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>29,-27,51,-27</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<connection>
<GID>9</GID>
<name>OUT_0</name></connection>
<intersection>38 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>38,-31.5,38,-27</points>
<connection>
<GID>7</GID>
<name>IN_0</name></connection>
<intersection>-27 1</intersection></vsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38,-43,38,-37.5</points>
<connection>
<GID>7</GID>
<name>OUT_0</name></connection>
<intersection>-43 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>38,-43,50.5,-43</points>
<connection>
<GID>3</GID>
<name>IN_1</name></connection>
<intersection>38 0</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47.5,-41,47.5,-29</points>
<intersection>-41 3</intersection>
<intersection>-35 2</intersection>
<intersection>-29 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47.5,-29,51,-29</points>
<connection>
<GID>2</GID>
<name>IN_1</name></connection>
<intersection>47.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>44.5,-35,47.5,-35</points>
<connection>
<GID>15</GID>
<name>OUT_0</name></connection>
<intersection>47.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>47.5,-41,50.5,-41</points>
<connection>
<GID>3</GID>
<name>IN_0</name></connection>
<intersection>47.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>57,-28,72,-28</points>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<connection>
<GID>2</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>64,-42,64,-40.5</points>
<intersection>-42 2</intersection>
<intersection>-40.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>64,-40.5,72,-40.5</points>
<connection>
<GID>5</GID>
<name>IN_1</name></connection>
<intersection>64 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>56.5,-42,64,-42</points>
<connection>
<GID>3</GID>
<name>OUT</name></connection>
<intersection>64 0</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>78,-39.5,91.5,-39.5</points>
<connection>
<GID>5</GID>
<name>OUT</name></connection>
<connection>
<GID>13</GID>
<name>N_in0</name></connection>
<intersection>79 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>79,-39.5,79,-30</points>
<intersection>-39.5 1</intersection>
<intersection>-30 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>72,-30,79,-30</points>
<connection>
<GID>4</GID>
<name>IN_1</name></connection>
<intersection>79 3</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>78,-29,92,-29</points>
<connection>
<GID>11</GID>
<name>N_in0</name></connection>
<connection>
<GID>4</GID>
<name>OUT</name></connection>
<intersection>81 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>81,-38.5,81,-29</points>
<intersection>-38.5 4</intersection>
<intersection>-29 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>72,-38.5,81,-38.5</points>
<connection>
<GID>5</GID>
<name>IN_0</name></connection>
<intersection>81 3</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-15.5,-70,47.5,-70</points>
<connection>
<GID>21</GID>
<name>IN_0</name></connection>
<intersection>-15.5 10</intersection>
<intersection>32.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>32.5,-74,32.5,-70</points>
<connection>
<GID>25</GID>
<name>IN_0</name></connection>
<intersection>-70 1</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>-15.5,-136,-15.5,-70</points>
<intersection>-136 11</intersection>
<intersection>-70 1</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>-37.5,-136,-15.5,-136</points>
<connection>
<GID>123</GID>
<name>OUT_0</name></connection>
<intersection>-15.5 10</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32.5,-83.5,32.5,-80</points>
<connection>
<GID>25</GID>
<name>OUT_0</name></connection>
<intersection>-83.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>32.5,-83.5,47,-83.5</points>
<connection>
<GID>22</GID>
<name>IN_1</name></connection>
<intersection>32.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>44,-81.5,44,-72</points>
<intersection>-81.5 3</intersection>
<intersection>-75 4</intersection>
<intersection>-72 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>44,-72,47.5,-72</points>
<connection>
<GID>21</GID>
<name>IN_1</name></connection>
<intersection>44 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>44,-81.5,47,-81.5</points>
<connection>
<GID>22</GID>
<name>IN_0</name></connection>
<intersection>44 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>42.5,-75,44,-75</points>
<connection>
<GID>35</GID>
<name>CLK</name></connection>
<intersection>44 0</intersection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53.5,-71,68.5,-71</points>
<connection>
<GID>21</GID>
<name>OUT</name></connection>
<connection>
<GID>23</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60.5,-82.5,60.5,-81</points>
<intersection>-82.5 2</intersection>
<intersection>-81 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>60.5,-81,68.5,-81</points>
<connection>
<GID>24</GID>
<name>IN_1</name></connection>
<intersection>60.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>53,-82.5,60.5,-82.5</points>
<connection>
<GID>22</GID>
<name>OUT</name></connection>
<intersection>60.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>74.5,-80,88,-80</points>
<connection>
<GID>24</GID>
<name>OUT</name></connection>
<connection>
<GID>28</GID>
<name>N_in0</name></connection>
<intersection>75.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>75.5,-80,75.5,-73</points>
<intersection>-80 1</intersection>
<intersection>-73 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>68.5,-73,75.5,-73</points>
<connection>
<GID>23</GID>
<name>IN_1</name></connection>
<intersection>75.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>74.5,-72,88.5,-72</points>
<connection>
<GID>23</GID>
<name>OUT</name></connection>
<connection>
<GID>27</GID>
<name>N_in0</name></connection>
<intersection>77.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>77.5,-79,77.5,-72</points>
<intersection>-79 4</intersection>
<intersection>-72 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>68.5,-79,77.5,-79</points>
<connection>
<GID>24</GID>
<name>IN_0</name></connection>
<intersection>77.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-25,-88,46,-88</points>
<connection>
<GID>36</GID>
<name>IN_0</name></connection>
<intersection>-25 6</intersection>
<intersection>31 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>31,-92,31,-88</points>
<connection>
<GID>40</GID>
<name>IN_0</name></connection>
<intersection>-88 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>-25,-134,-25,-88</points>
<intersection>-134 7</intersection>
<intersection>-88 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-37.5,-134,-25,-134</points>
<connection>
<GID>123</GID>
<name>OUT_1</name></connection>
<intersection>-25 6</intersection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31,-104,31,-98</points>
<connection>
<GID>40</GID>
<name>OUT_0</name></connection>
<intersection>-104 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>31,-104,45.5,-104</points>
<connection>
<GID>37</GID>
<name>IN_1</name></connection>
<intersection>31 0</intersection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>42.5,-102,42.5,-90</points>
<intersection>-102 3</intersection>
<intersection>-95.5 4</intersection>
<intersection>-90 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>42.5,-90,46,-90</points>
<connection>
<GID>36</GID>
<name>IN_1</name></connection>
<intersection>42.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>42.5,-102,45.5,-102</points>
<connection>
<GID>37</GID>
<name>IN_0</name></connection>
<intersection>42.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>41,-95.5,42.5,-95.5</points>
<connection>
<GID>47</GID>
<name>CLK</name></connection>
<intersection>42.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>52,-89,67,-89</points>
<connection>
<GID>38</GID>
<name>IN_0</name></connection>
<connection>
<GID>36</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>59,-103,59,-101.5</points>
<intersection>-103 2</intersection>
<intersection>-101.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>59,-101.5,67,-101.5</points>
<connection>
<GID>39</GID>
<name>IN_1</name></connection>
<intersection>59 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>51.5,-103,59,-103</points>
<connection>
<GID>37</GID>
<name>OUT</name></connection>
<intersection>59 0</intersection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73,-100.5,86.5,-100.5</points>
<connection>
<GID>39</GID>
<name>OUT</name></connection>
<connection>
<GID>43</GID>
<name>N_in0</name></connection>
<intersection>74 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>74,-100.5,74,-91</points>
<intersection>-100.5 1</intersection>
<intersection>-91 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>67,-91,74,-91</points>
<connection>
<GID>38</GID>
<name>IN_1</name></connection>
<intersection>74 3</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73,-90,87,-90</points>
<connection>
<GID>42</GID>
<name>N_in0</name></connection>
<connection>
<GID>38</GID>
<name>OUT</name></connection>
<intersection>76 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>76,-99.5,76,-90</points>
<intersection>-99.5 4</intersection>
<intersection>-90 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>67,-99.5,76,-99.5</points>
<connection>
<GID>39</GID>
<name>IN_0</name></connection>
<intersection>76 3</intersection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-30,-110,46.5,-110</points>
<connection>
<GID>48</GID>
<name>IN_0</name></connection>
<intersection>-30 6</intersection>
<intersection>31.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>31.5,-114,31.5,-110</points>
<connection>
<GID>52</GID>
<name>IN_0</name></connection>
<intersection>-110 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>-30,-132,-30,-110</points>
<intersection>-132 7</intersection>
<intersection>-110 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-37.5,-132,-30,-132</points>
<connection>
<GID>123</GID>
<name>OUT_2</name></connection>
<intersection>-30 6</intersection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31.5,-126,31.5,-120</points>
<connection>
<GID>52</GID>
<name>OUT_0</name></connection>
<intersection>-126 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>31.5,-126,46,-126</points>
<connection>
<GID>49</GID>
<name>IN_1</name></connection>
<intersection>31.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43,-124,43,-112</points>
<intersection>-124 3</intersection>
<intersection>-117.5 4</intersection>
<intersection>-112 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>43,-112,46.5,-112</points>
<connection>
<GID>48</GID>
<name>IN_1</name></connection>
<intersection>43 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>43,-124,46,-124</points>
<connection>
<GID>49</GID>
<name>IN_0</name></connection>
<intersection>43 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>41.5,-117.5,43,-117.5</points>
<connection>
<GID>59</GID>
<name>CLK</name></connection>
<intersection>43 0</intersection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>52.5,-111,67.5,-111</points>
<connection>
<GID>50</GID>
<name>IN_0</name></connection>
<connection>
<GID>48</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>59.5,-125,59.5,-123.5</points>
<intersection>-125 2</intersection>
<intersection>-123.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>59.5,-123.5,67.5,-123.5</points>
<connection>
<GID>51</GID>
<name>IN_1</name></connection>
<intersection>59.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>52,-125,59.5,-125</points>
<connection>
<GID>49</GID>
<name>OUT</name></connection>
<intersection>59.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73.5,-122.5,87,-122.5</points>
<connection>
<GID>55</GID>
<name>N_in0</name></connection>
<connection>
<GID>51</GID>
<name>OUT</name></connection>
<intersection>74.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>74.5,-122.5,74.5,-113</points>
<intersection>-122.5 1</intersection>
<intersection>-113 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>67.5,-113,74.5,-113</points>
<connection>
<GID>50</GID>
<name>IN_1</name></connection>
<intersection>74.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73.5,-112,87.5,-112</points>
<connection>
<GID>54</GID>
<name>N_in0</name></connection>
<connection>
<GID>50</GID>
<name>OUT</name></connection>
<intersection>76.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>76.5,-121.5,76.5,-112</points>
<intersection>-121.5 4</intersection>
<intersection>-112 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>67.5,-121.5,76.5,-121.5</points>
<connection>
<GID>51</GID>
<name>IN_0</name></connection>
<intersection>76.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-37.5,-130.5,47.5,-130.5</points>
<intersection>-37.5 6</intersection>
<intersection>32.5 3</intersection>
<intersection>47.5 8</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>32.5,-136.5,32.5,-130.5</points>
<connection>
<GID>64</GID>
<name>IN_0</name></connection>
<intersection>-130.5 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>-37.5,-130.5,-37.5,-130</points>
<connection>
<GID>123</GID>
<name>OUT_3</name></connection>
<intersection>-130.5 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>47.5,-132.5,47.5,-130.5</points>
<connection>
<GID>60</GID>
<name>IN_0</name></connection>
<intersection>-130.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32.5,-148.5,32.5,-142.5</points>
<connection>
<GID>64</GID>
<name>OUT_0</name></connection>
<intersection>-148.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>32.5,-148.5,47,-148.5</points>
<connection>
<GID>61</GID>
<name>IN_1</name></connection>
<intersection>32.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>44,-146.5,44,-134.5</points>
<intersection>-146.5 3</intersection>
<intersection>-140 4</intersection>
<intersection>-134.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>44,-134.5,47.5,-134.5</points>
<connection>
<GID>60</GID>
<name>IN_1</name></connection>
<intersection>44 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>44,-146.5,47,-146.5</points>
<connection>
<GID>61</GID>
<name>IN_0</name></connection>
<intersection>44 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>42.5,-140,44,-140</points>
<connection>
<GID>71</GID>
<name>CLK</name></connection>
<intersection>44 0</intersection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53.5,-133.5,68.5,-133.5</points>
<connection>
<GID>62</GID>
<name>IN_0</name></connection>
<connection>
<GID>60</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60.5,-147.5,60.5,-146</points>
<intersection>-147.5 2</intersection>
<intersection>-146 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>60.5,-146,68.5,-146</points>
<connection>
<GID>63</GID>
<name>IN_1</name></connection>
<intersection>60.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>53,-147.5,60.5,-147.5</points>
<connection>
<GID>61</GID>
<name>OUT</name></connection>
<intersection>60.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>74.5,-145,88,-145</points>
<connection>
<GID>67</GID>
<name>N_in0</name></connection>
<connection>
<GID>63</GID>
<name>OUT</name></connection>
<intersection>75.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>75.5,-145,75.5,-135.5</points>
<intersection>-145 1</intersection>
<intersection>-135.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>68.5,-135.5,75.5,-135.5</points>
<connection>
<GID>62</GID>
<name>IN_1</name></connection>
<intersection>75.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>74.5,-134.5,88.5,-134.5</points>
<connection>
<GID>66</GID>
<name>N_in0</name></connection>
<connection>
<GID>62</GID>
<name>OUT</name></connection>
<intersection>77.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>77.5,-144,77.5,-134.5</points>
<intersection>-144 4</intersection>
<intersection>-134.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>68.5,-144,77.5,-144</points>
<connection>
<GID>63</GID>
<name>IN_0</name></connection>
<intersection>77.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>71</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-15.5,-157.5,47.5,-157.5</points>
<connection>
<GID>136</GID>
<name>IN_0</name></connection>
<intersection>-15.5 10</intersection>
<intersection>32.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>32.5,-161.5,32.5,-157.5</points>
<connection>
<GID>140</GID>
<name>IN_0</name></connection>
<intersection>-157.5 1</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>-15.5,-157.5,-15.5,-155</points>
<intersection>-157.5 1</intersection>
<intersection>-155 11</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>-38,-155,-15.5,-155</points>
<connection>
<GID>176</GID>
<name>OUT_0</name></connection>
<intersection>-15.5 10</intersection></hsegment></shape></wire>
<wire>
<ID>72</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32.5,-171,32.5,-167.5</points>
<connection>
<GID>140</GID>
<name>OUT_0</name></connection>
<intersection>-171 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>32.5,-171,47,-171</points>
<connection>
<GID>137</GID>
<name>IN_1</name></connection>
<intersection>32.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>73</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>44,-169,44,-159.5</points>
<intersection>-169 3</intersection>
<intersection>-162.5 4</intersection>
<intersection>-159.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>44,-159.5,47.5,-159.5</points>
<connection>
<GID>136</GID>
<name>IN_1</name></connection>
<intersection>44 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>44,-169,47,-169</points>
<connection>
<GID>137</GID>
<name>IN_0</name></connection>
<intersection>44 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>42.5,-162.5,44,-162.5</points>
<connection>
<GID>145</GID>
<name>CLK</name></connection>
<intersection>44 0</intersection></hsegment></shape></wire>
<wire>
<ID>74</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53.5,-158.5,68.5,-158.5</points>
<connection>
<GID>136</GID>
<name>OUT</name></connection>
<connection>
<GID>138</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>75</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60.5,-170,60.5,-168.5</points>
<intersection>-170 2</intersection>
<intersection>-168.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>60.5,-168.5,68.5,-168.5</points>
<connection>
<GID>139</GID>
<name>IN_1</name></connection>
<intersection>60.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>53,-170,60.5,-170</points>
<connection>
<GID>137</GID>
<name>OUT</name></connection>
<intersection>60.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>76</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>74.5,-167.5,88,-167.5</points>
<connection>
<GID>139</GID>
<name>OUT</name></connection>
<connection>
<GID>142</GID>
<name>N_in0</name></connection>
<intersection>75.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>75.5,-167.5,75.5,-160.5</points>
<intersection>-167.5 1</intersection>
<intersection>-160.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>68.5,-160.5,75.5,-160.5</points>
<connection>
<GID>138</GID>
<name>IN_1</name></connection>
<intersection>75.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>77</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>74.5,-159.5,88.5,-159.5</points>
<connection>
<GID>138</GID>
<name>OUT</name></connection>
<connection>
<GID>141</GID>
<name>N_in0</name></connection>
<intersection>77.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>77.5,-166.5,77.5,-159.5</points>
<intersection>-166.5 4</intersection>
<intersection>-159.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>68.5,-166.5,77.5,-166.5</points>
<connection>
<GID>139</GID>
<name>IN_0</name></connection>
<intersection>77.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>78</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-25,-175.5,46,-175.5</points>
<connection>
<GID>146</GID>
<name>IN_0</name></connection>
<intersection>-25 6</intersection>
<intersection>31 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>31,-179.5,31,-175.5</points>
<connection>
<GID>150</GID>
<name>IN_0</name></connection>
<intersection>-175.5 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>-25,-175.5,-25,-153</points>
<intersection>-175.5 1</intersection>
<intersection>-153 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-38,-153,-25,-153</points>
<connection>
<GID>176</GID>
<name>OUT_1</name></connection>
<intersection>-25 6</intersection></hsegment></shape></wire>
<wire>
<ID>79</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31,-191.5,31,-185.5</points>
<connection>
<GID>150</GID>
<name>OUT_0</name></connection>
<intersection>-191.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>31,-191.5,45.5,-191.5</points>
<connection>
<GID>147</GID>
<name>IN_1</name></connection>
<intersection>31 0</intersection></hsegment></shape></wire>
<wire>
<ID>80</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>42.5,-189.5,42.5,-177.5</points>
<intersection>-189.5 3</intersection>
<intersection>-183 4</intersection>
<intersection>-177.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>42.5,-177.5,46,-177.5</points>
<connection>
<GID>146</GID>
<name>IN_1</name></connection>
<intersection>42.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>42.5,-189.5,45.5,-189.5</points>
<connection>
<GID>147</GID>
<name>IN_0</name></connection>
<intersection>42.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>41,-183,42.5,-183</points>
<connection>
<GID>155</GID>
<name>CLK</name></connection>
<intersection>42.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>81</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>52,-176.5,67,-176.5</points>
<connection>
<GID>146</GID>
<name>OUT</name></connection>
<connection>
<GID>148</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>82</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>59,-190.5,59,-189</points>
<intersection>-190.5 2</intersection>
<intersection>-189 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>59,-189,67,-189</points>
<connection>
<GID>149</GID>
<name>IN_1</name></connection>
<intersection>59 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>51.5,-190.5,59,-190.5</points>
<connection>
<GID>147</GID>
<name>OUT</name></connection>
<intersection>59 0</intersection></hsegment></shape></wire>
<wire>
<ID>83</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73,-188,86.5,-188</points>
<connection>
<GID>149</GID>
<name>OUT</name></connection>
<connection>
<GID>152</GID>
<name>N_in0</name></connection>
<intersection>74 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>74,-188,74,-178.5</points>
<intersection>-188 1</intersection>
<intersection>-178.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>67,-178.5,74,-178.5</points>
<connection>
<GID>148</GID>
<name>IN_1</name></connection>
<intersection>74 3</intersection></hsegment></shape></wire>
<wire>
<ID>84</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73,-177.5,87,-177.5</points>
<connection>
<GID>148</GID>
<name>OUT</name></connection>
<connection>
<GID>151</GID>
<name>N_in0</name></connection>
<intersection>76 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>76,-187,76,-177.5</points>
<intersection>-187 4</intersection>
<intersection>-177.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>67,-187,76,-187</points>
<connection>
<GID>149</GID>
<name>IN_0</name></connection>
<intersection>76 3</intersection></hsegment></shape></wire>
<wire>
<ID>85</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-30,-197.5,46.5,-197.5</points>
<connection>
<GID>156</GID>
<name>IN_0</name></connection>
<intersection>-30 6</intersection>
<intersection>31.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>31.5,-201.5,31.5,-197.5</points>
<connection>
<GID>160</GID>
<name>IN_0</name></connection>
<intersection>-197.5 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>-30,-197.5,-30,-151</points>
<intersection>-197.5 1</intersection>
<intersection>-151 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-38,-151,-30,-151</points>
<connection>
<GID>176</GID>
<name>OUT_2</name></connection>
<intersection>-30 6</intersection></hsegment></shape></wire>
<wire>
<ID>86</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31.5,-213.5,31.5,-207.5</points>
<connection>
<GID>160</GID>
<name>OUT_0</name></connection>
<intersection>-213.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>31.5,-213.5,46,-213.5</points>
<connection>
<GID>157</GID>
<name>IN_1</name></connection>
<intersection>31.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>87</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43,-211.5,43,-199.5</points>
<intersection>-211.5 3</intersection>
<intersection>-205 4</intersection>
<intersection>-199.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>43,-199.5,46.5,-199.5</points>
<connection>
<GID>156</GID>
<name>IN_1</name></connection>
<intersection>43 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>43,-211.5,46,-211.5</points>
<connection>
<GID>157</GID>
<name>IN_0</name></connection>
<intersection>43 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>41.5,-205,43,-205</points>
<connection>
<GID>165</GID>
<name>CLK</name></connection>
<intersection>43 0</intersection></hsegment></shape></wire>
<wire>
<ID>88</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>52.5,-198.5,67.5,-198.5</points>
<connection>
<GID>156</GID>
<name>OUT</name></connection>
<connection>
<GID>158</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>89</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>59.5,-212.5,59.5,-211</points>
<intersection>-212.5 2</intersection>
<intersection>-211 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>59.5,-211,67.5,-211</points>
<connection>
<GID>159</GID>
<name>IN_1</name></connection>
<intersection>59.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>52,-212.5,59.5,-212.5</points>
<connection>
<GID>157</GID>
<name>OUT</name></connection>
<intersection>59.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>90</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73.5,-210,87,-210</points>
<connection>
<GID>159</GID>
<name>OUT</name></connection>
<connection>
<GID>162</GID>
<name>N_in0</name></connection>
<intersection>74.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>74.5,-210,74.5,-200.5</points>
<intersection>-210 1</intersection>
<intersection>-200.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>67.5,-200.5,74.5,-200.5</points>
<connection>
<GID>158</GID>
<name>IN_1</name></connection>
<intersection>74.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>91</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73.5,-199.5,87.5,-199.5</points>
<connection>
<GID>158</GID>
<name>OUT</name></connection>
<connection>
<GID>161</GID>
<name>N_in0</name></connection>
<intersection>76.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>76.5,-209,76.5,-199.5</points>
<intersection>-209 4</intersection>
<intersection>-199.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>67.5,-209,76.5,-209</points>
<connection>
<GID>159</GID>
<name>IN_0</name></connection>
<intersection>76.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>92</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-37.5,-218,47.5,-218</points>
<intersection>-37.5 6</intersection>
<intersection>32.5 3</intersection>
<intersection>47.5 8</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>32.5,-224,32.5,-218</points>
<connection>
<GID>170</GID>
<name>IN_0</name></connection>
<intersection>-218 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>-37.5,-218,-37.5,-149</points>
<intersection>-218 1</intersection>
<intersection>-149 15</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>47.5,-220,47.5,-218</points>
<connection>
<GID>166</GID>
<name>IN_0</name></connection>
<intersection>-218 1</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>-38,-149,-37.5,-149</points>
<connection>
<GID>176</GID>
<name>OUT_3</name></connection>
<intersection>-37.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>93</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32.5,-236,32.5,-230</points>
<connection>
<GID>170</GID>
<name>OUT_0</name></connection>
<intersection>-236 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>32.5,-236,47,-236</points>
<connection>
<GID>167</GID>
<name>IN_1</name></connection>
<intersection>32.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>94</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>44,-234,44,-222</points>
<intersection>-234 3</intersection>
<intersection>-227.5 4</intersection>
<intersection>-222 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>44,-222,47.5,-222</points>
<connection>
<GID>166</GID>
<name>IN_1</name></connection>
<intersection>44 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>44,-234,47,-234</points>
<connection>
<GID>167</GID>
<name>IN_0</name></connection>
<intersection>44 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>42.5,-227.5,44,-227.5</points>
<connection>
<GID>175</GID>
<name>CLK</name></connection>
<intersection>44 0</intersection></hsegment></shape></wire>
<wire>
<ID>95</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53.5,-221,68.5,-221</points>
<connection>
<GID>166</GID>
<name>OUT</name></connection>
<connection>
<GID>168</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>96</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60.5,-235,60.5,-233.5</points>
<intersection>-235 2</intersection>
<intersection>-233.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>60.5,-233.5,68.5,-233.5</points>
<connection>
<GID>169</GID>
<name>IN_1</name></connection>
<intersection>60.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>53,-235,60.5,-235</points>
<connection>
<GID>167</GID>
<name>OUT</name></connection>
<intersection>60.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>97</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>74.5,-232.5,88,-232.5</points>
<connection>
<GID>169</GID>
<name>OUT</name></connection>
<connection>
<GID>172</GID>
<name>N_in0</name></connection>
<intersection>75.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>75.5,-232.5,75.5,-223</points>
<intersection>-232.5 1</intersection>
<intersection>-223 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>68.5,-223,75.5,-223</points>
<connection>
<GID>168</GID>
<name>IN_1</name></connection>
<intersection>75.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>98</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>74.5,-222,88.5,-222</points>
<connection>
<GID>168</GID>
<name>OUT</name></connection>
<connection>
<GID>171</GID>
<name>N_in0</name></connection>
<intersection>77.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>77.5,-231.5,77.5,-222</points>
<intersection>-231.5 4</intersection>
<intersection>-222 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>68.5,-231.5,77.5,-231.5</points>
<connection>
<GID>169</GID>
<name>IN_0</name></connection>
<intersection>77.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>99</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>123.5,-147,123.5,-72</points>
<intersection>-147 1</intersection>
<intersection>-72 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>123.5,-147,159,-147</points>
<connection>
<GID>178</GID>
<name>IN_0</name></connection>
<intersection>123.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>90.5,-72,123.5,-72</points>
<connection>
<GID>27</GID>
<name>N_in1</name></connection>
<intersection>123.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>100</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>122.5,-146,122.5,-90</points>
<intersection>-146 1</intersection>
<intersection>-90 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>122.5,-146,159,-146</points>
<connection>
<GID>178</GID>
<name>IN_1</name></connection>
<intersection>122.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>89,-90,122.5,-90</points>
<connection>
<GID>42</GID>
<name>N_in1</name></connection>
<intersection>122.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>101</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>123,-145,123,-112</points>
<intersection>-145 1</intersection>
<intersection>-112 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>123,-145,159,-145</points>
<connection>
<GID>178</GID>
<name>IN_2</name></connection>
<intersection>123 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>89.5,-112,123,-112</points>
<connection>
<GID>54</GID>
<name>N_in1</name></connection>
<intersection>123 0</intersection></hsegment></shape></wire>
<wire>
<ID>102</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>123.5,-144,123.5,-134.5</points>
<intersection>-144 1</intersection>
<intersection>-134.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>123.5,-144,159,-144</points>
<connection>
<GID>178</GID>
<name>IN_3</name></connection>
<intersection>123.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>90.5,-134.5,123.5,-134.5</points>
<connection>
<GID>66</GID>
<name>N_in1</name></connection>
<intersection>123.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>103</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>123.5,-159.5,123.5,-143</points>
<intersection>-159.5 2</intersection>
<intersection>-143 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>123.5,-143,159,-143</points>
<connection>
<GID>178</GID>
<name>IN_4</name></connection>
<intersection>123.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>90.5,-159.5,123.5,-159.5</points>
<connection>
<GID>141</GID>
<name>N_in1</name></connection>
<intersection>123.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>104</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>123,-177.5,123,-142</points>
<intersection>-177.5 2</intersection>
<intersection>-142 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>123,-142,159,-142</points>
<connection>
<GID>178</GID>
<name>IN_5</name></connection>
<intersection>123 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>89,-177.5,123,-177.5</points>
<connection>
<GID>151</GID>
<name>N_in1</name></connection>
<intersection>123 0</intersection></hsegment></shape></wire>
<wire>
<ID>105</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>123,-199.5,123,-141</points>
<intersection>-199.5 2</intersection>
<intersection>-141 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>123,-141,159,-141</points>
<connection>
<GID>178</GID>
<name>IN_6</name></connection>
<intersection>123 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>89.5,-199.5,123,-199.5</points>
<connection>
<GID>161</GID>
<name>N_in1</name></connection>
<intersection>123 0</intersection></hsegment></shape></wire>
<wire>
<ID>106</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>123.5,-222,123.5,-140</points>
<intersection>-222 2</intersection>
<intersection>-140 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>123.5,-140,159,-140</points>
<connection>
<GID>178</GID>
<name>IN_7</name></connection>
<intersection>123.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>90.5,-222,123.5,-222</points>
<connection>
<GID>171</GID>
<name>N_in1</name></connection>
<intersection>123.5 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,0,177.8,-91.7</PageViewport></page 1>
<page 2>
<PageViewport>0,0,177.8,-91.7</PageViewport></page 2>
<page 3>
<PageViewport>0,0,177.8,-91.7</PageViewport></page 3>
<page 4>
<PageViewport>0,0,177.8,-91.7</PageViewport></page 4>
<page 5>
<PageViewport>0,0,177.8,-91.7</PageViewport></page 5>
<page 6>
<PageViewport>0,0,177.8,-91.7</PageViewport></page 6>
<page 7>
<PageViewport>0,0,177.8,-91.7</PageViewport></page 7>
<page 8>
<PageViewport>0,0,177.8,-91.7</PageViewport></page 8>
<page 9>
<PageViewport>0,0,177.8,-91.7</PageViewport></page 9></circuit>